library ieee;
use ieee.std_logic_1164.all;

entity Sin_Gen_Peripheral is
port(
	CPU_reset:	in	std_logic;
	CPU_clk:	in	std_logic;
	clk_50:		in	std_logic;
	
	En_Amp1:		in	std_logic;
	input_Amp1:		in	std_logic_vector(13 downto 0);
	output_Amp1:	out	std_logic_vector(13 downto 0);
	
	En_Amp2:		in	std_logic;
	input_Amp2:		in	std_logic_vector(13 downto 0);
	output_Amp2:	out	std_logic_vector(13 downto 0);
	
	En_phase1:		in	std_logic;
	input_phase1:	in	std_logic_vector(12 downto 0);
	output_phase1:	out	std_logic_vector(12 downto 0);
	
	En_phase2:		in	std_logic;
	input_phase2:	in	std_logic_vector(12 downto 0);
	output_phase2:	out	std_logic_vector(12 downto 0);
	
	DAC_MODE:		out	std_logic;
	DAC_WRT_A:		out	std_logic;
	DAC_WRT_B:		out	std_logic;
	DAC_CLK_A:		out	std_logic;
	DAC_CLK_B:		out	std_logic;
	DAC_DA:			out	std_logic_vector(13 downto 0);
	DAC_DB:			out	std_logic_vector(13 downto 0));
end;

architecture one of Sin_Gen_Peripheral is
	
	-- / Components \ --
	component sin_Gen
	port(
		reset:		in	std_logic;
		clk:		in	std_logic;
		amplitude1:	in	std_logic_vector(13 downto 0);
		phase_inc1:	in	std_logic_vector(12 downto 0);
		amplitude2:	in	std_logic_vector(13 downto 0);
		phase_inc2:	in	std_logic_vector(12 downto 0);
		outpt:		out	std_logic_vector(13 downto 0));
	end component;
	
	component PLL
	port(
		areset:	in	std_logic;
		inclk0:	in	std_logic;
		c0:		out	std_logic);
	end component;

	component sin_Gen_Peripheral_Register
	generic(Bits:integer:=32);
	port(
		reset:	in	std_logic;
		clk:	in	std_logic;
		En:		in	std_logic;
		input:	in	std_logic_vector(Bits-1 downto 0);
		output:	out	std_logic_vector(Bits-1 downto 0));
	end component;
	-- / Components \ --
	
	-- / Signals \ --
	signal clk_125:			std_logic;
	signal sig_output_Amp1:	std_logic_vector(13 downto 0);
	signal sig_output_Amp2:	std_logic_vector(13 downto 0);
	signal sig_output_phase1:	std_logic_vector(12 downto 0);
	signal sig_output_phase2:	std_logic_vector(12 downto 0);
	signal sin_signal:			std_logic_vector(13 downto 0);
	-- / Signals \ --
	
begin
	
	U1: PLL port map(
		areset	=>	'0',
		inclk0	=>	clk_50,		--	50[MHz]  clk signal input
		c0		=>	clk_125);	--	125[MHz] clk signal output
	
	U2: sin_Gen port map(
		reset	=>	CPU_reset,
		clk		=>	clk_125,
		
		amplitude1	=>	sig_output_Amp1,
		phase_inc1	=>	sig_output_phase1,
		amplitude2	=>	sig_output_Amp2,
		phase_inc2	=>	sig_output_phase2,
		
		outpt		=>	sin_signal);
	
	Amp1:	sin_Gen_Peripheral_Register generic map(14) port map(
		reset	=>	CPU_reset,
		clk		=>	CPU_clk,
		En		=>	En_Amp1,
		input	=>	input_Amp1,
		output	=>	sig_output_Amp1);
	output_Amp1 <= sig_output_Amp1;
	
	Amp2:	sin_Gen_Peripheral_Register generic map(14) port map(
		reset	=>	CPU_reset,
		clk		=>	CPU_clk,
		En		=>	En_Amp2,
		input	=>	input_Amp2,
		output	=>	sig_output_Amp2);
	output_Amp2 <= sig_output_Amp2;
	
	phase1:	sin_Gen_Peripheral_Register generic map(13) port map(
		reset	=>	CPU_reset,
		clk		=>	CPU_clk,
		En		=>	En_phase1,
		input	=>	input_phase1,
		output	=>	sig_output_phase1);
	output_phase1 <= sig_output_phase1;
	
	phase2:	sin_Gen_Peripheral_Register generic map(13) port map(
		reset	=>	CPU_reset,
		clk		=>	CPU_clk,
		En		=>	En_phase2,
		input	=>	input_phase2,
		output	=>	sig_output_phase2);
	output_phase2 <= sig_output_phase2;
	
	DAC_MODE <= '1';
	
	DAC_WRT_A <= clk_125;
	DAC_WRT_B <= clk_125;
	
	DAC_CLK_A <= clk_125;
	DAC_CLK_B <= clk_125;
	
	DAC_DA <= (not sin_signal(13)) & sin_signal(12 downto 0);
	
	DAC_DB <= (not sin_signal(13)) & sin_signal(12 downto 0);
	
end;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;

entity sin_Gen is
port(
	reset:	in		std_logic;
	clk:		in		std_logic;
	
	amplitude1:	in	std_logic_vector(13 downto 0);
	phase_inc1:	in	std_logic_vector(12 downto 0);
	amplitude2:	in	std_logic_vector(13 downto 0);
	phase_inc2:	in	std_logic_vector(12 downto 0);
	
	outpt:	out	std_logic_vector(13 downto 0));
end;

architecture one of sin_Gen is
	-- / Components \ --
	component sin_rom
	port(
		address1:	in		std_logic_vector(12 downto 0);
		amplitude1:	in		std_logic_vector(13 downto 0);
		data_out1:	out	std_logic_vector(13 downto 0);
		
		address2:	in		std_logic_vector(12 downto 0);
		amplitude2:	in		std_logic_vector(13 downto 0);
		data_out2:	out	std_logic_vector(13 downto 0));
	end component;
	
	component sin_counter
	port(
		reset:	in		std_logic;
		clk:		in		std_logic;
		phase_inc:	in	std_logic_vector(12 downto 0);
		Q:			out	std_logic_vector(12 downto 0));
	end component;
	-- / Components \ --
	
	-- / Signals \ --
	signal Q1:			std_logic_vector(12 downto 0);
	signal Q2:			std_logic_vector(12 downto 0);
	
	signal outpt1:		std_logic_vector(13 downto 0);
	signal outpt2:		std_logic_vector(13 downto 0);
	-- / Signals \ --
begin
	
	U1:	sin_counter port map(
		reset			=>	reset,
		clk			=>	clk,
		phase_inc	=> phase_inc1,
		Q				=>	Q1);
	
	U2:	sin_counter port map(
		reset			=>	reset,
		clk			=>	clk,
		phase_inc	=> phase_inc2,
		Q				=>	Q2);
	
	U3:	sin_rom port map(
		address1		=>	Q1,
		amplitude1	=>	amplitude1,
		data_out1	=>	outpt1,
		
		address2		=>	Q2,
		amplitude2	=>	amplitude2,
		data_out2	=>	outpt2);
		
		outpt <= outpt1 + outpt2;
end;

-- SubModule: sin_rom --

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use ieee.std_logic_arith.all;

entity sin_rom is
port(
	address1:	in		std_logic_vector(12 downto 0);
	amplitude1:	in		std_logic_vector(13 downto 0);	-- 14[Bits], 12[Bits] fraction
	data_out1:	out	std_logic_vector(13 downto 0);
	
	address2:	in		std_logic_vector(12 downto 0);
	amplitude2:	in		std_logic_vector(13 downto 0);
	data_out2:	out	std_logic_vector(13 downto 0));
end;

architecture one of sin_rom is
	
	type lut_rom is array(-4096 to 4095) of std_logic_vector(13 downto 0);
	signal rom:lut_rom:=
	(	conv_std_logic_vector(0,14),
		conv_std_logic_vector(6,14),
		conv_std_logic_vector(12,14),
		conv_std_logic_vector(18,14),
		conv_std_logic_vector(25,14),
		conv_std_logic_vector(31,14),
		conv_std_logic_vector(37,14),
		conv_std_logic_vector(43,14),
		conv_std_logic_vector(50,14),
		conv_std_logic_vector(56,14),
		conv_std_logic_vector(62,14),
		conv_std_logic_vector(69,14),
		conv_std_logic_vector(75,14),
		conv_std_logic_vector(81,14),
		conv_std_logic_vector(87,14),
		conv_std_logic_vector(94,14),
		conv_std_logic_vector(100,14),
		conv_std_logic_vector(106,14),
		conv_std_logic_vector(113,14),
		conv_std_logic_vector(119,14),
		conv_std_logic_vector(125,14),
		conv_std_logic_vector(131,14),
		conv_std_logic_vector(138,14),
		conv_std_logic_vector(144,14),
		conv_std_logic_vector(150,14),
		conv_std_logic_vector(157,14),
		conv_std_logic_vector(163,14),
		conv_std_logic_vector(169,14),
		conv_std_logic_vector(175,14),
		conv_std_logic_vector(182,14),
		conv_std_logic_vector(188,14),
		conv_std_logic_vector(194,14),
		conv_std_logic_vector(201,14),
		conv_std_logic_vector(207,14),
		conv_std_logic_vector(213,14),
		conv_std_logic_vector(219,14),
		conv_std_logic_vector(226,14),
		conv_std_logic_vector(232,14),
		conv_std_logic_vector(238,14),
		conv_std_logic_vector(245,14),
		conv_std_logic_vector(251,14),
		conv_std_logic_vector(257,14),
		conv_std_logic_vector(263,14),
		conv_std_logic_vector(270,14),
		conv_std_logic_vector(276,14),
		conv_std_logic_vector(282,14),
		conv_std_logic_vector(288,14),
		conv_std_logic_vector(295,14),
		conv_std_logic_vector(301,14),
		conv_std_logic_vector(307,14),
		conv_std_logic_vector(314,14),
		conv_std_logic_vector(320,14),
		conv_std_logic_vector(326,14),
		conv_std_logic_vector(332,14),
		conv_std_logic_vector(339,14),
		conv_std_logic_vector(345,14),
		conv_std_logic_vector(351,14),
		conv_std_logic_vector(358,14),
		conv_std_logic_vector(364,14),
		conv_std_logic_vector(370,14),
		conv_std_logic_vector(376,14),
		conv_std_logic_vector(383,14),
		conv_std_logic_vector(389,14),
		conv_std_logic_vector(395,14),
		conv_std_logic_vector(401,14),
		conv_std_logic_vector(408,14),
		conv_std_logic_vector(414,14),
		conv_std_logic_vector(420,14),
		conv_std_logic_vector(427,14),
		conv_std_logic_vector(433,14),
		conv_std_logic_vector(439,14),
		conv_std_logic_vector(445,14),
		conv_std_logic_vector(452,14),
		conv_std_logic_vector(458,14),
		conv_std_logic_vector(464,14),
		conv_std_logic_vector(470,14),
		conv_std_logic_vector(477,14),
		conv_std_logic_vector(483,14),
		conv_std_logic_vector(489,14),
		conv_std_logic_vector(496,14),
		conv_std_logic_vector(502,14),
		conv_std_logic_vector(508,14),
		conv_std_logic_vector(514,14),
		conv_std_logic_vector(521,14),
		conv_std_logic_vector(527,14),
		conv_std_logic_vector(533,14),
		conv_std_logic_vector(539,14),
		conv_std_logic_vector(546,14),
		conv_std_logic_vector(552,14),
		conv_std_logic_vector(558,14),
		conv_std_logic_vector(565,14),
		conv_std_logic_vector(571,14),
		conv_std_logic_vector(577,14),
		conv_std_logic_vector(583,14),
		conv_std_logic_vector(590,14),
		conv_std_logic_vector(596,14),
		conv_std_logic_vector(602,14),
		conv_std_logic_vector(608,14),
		conv_std_logic_vector(615,14),
		conv_std_logic_vector(621,14),
		conv_std_logic_vector(627,14),
		conv_std_logic_vector(633,14),
		conv_std_logic_vector(640,14),
		conv_std_logic_vector(646,14),
		conv_std_logic_vector(652,14),
		conv_std_logic_vector(659,14),
		conv_std_logic_vector(665,14),
		conv_std_logic_vector(671,14),
		conv_std_logic_vector(677,14),
		conv_std_logic_vector(684,14),
		conv_std_logic_vector(690,14),
		conv_std_logic_vector(696,14),
		conv_std_logic_vector(702,14),
		conv_std_logic_vector(709,14),
		conv_std_logic_vector(715,14),
		conv_std_logic_vector(721,14),
		conv_std_logic_vector(727,14),
		conv_std_logic_vector(734,14),
		conv_std_logic_vector(740,14),
		conv_std_logic_vector(746,14),
		conv_std_logic_vector(752,14),
		conv_std_logic_vector(759,14),
		conv_std_logic_vector(765,14),
		conv_std_logic_vector(771,14),
		conv_std_logic_vector(777,14),
		conv_std_logic_vector(784,14),
		conv_std_logic_vector(790,14),
		conv_std_logic_vector(796,14),
		conv_std_logic_vector(802,14),
		conv_std_logic_vector(809,14),
		conv_std_logic_vector(815,14),
		conv_std_logic_vector(821,14),
		conv_std_logic_vector(827,14),
		conv_std_logic_vector(834,14),
		conv_std_logic_vector(840,14),
		conv_std_logic_vector(846,14),
		conv_std_logic_vector(852,14),
		conv_std_logic_vector(859,14),
		conv_std_logic_vector(865,14),
		conv_std_logic_vector(871,14),
		conv_std_logic_vector(877,14),
		conv_std_logic_vector(884,14),
		conv_std_logic_vector(890,14),
		conv_std_logic_vector(896,14),
		conv_std_logic_vector(902,14),
		conv_std_logic_vector(909,14),
		conv_std_logic_vector(915,14),
		conv_std_logic_vector(921,14),
		conv_std_logic_vector(927,14),
		conv_std_logic_vector(934,14),
		conv_std_logic_vector(940,14),
		conv_std_logic_vector(946,14),
		conv_std_logic_vector(952,14),
		conv_std_logic_vector(959,14),
		conv_std_logic_vector(965,14),
		conv_std_logic_vector(971,14),
		conv_std_logic_vector(977,14),
		conv_std_logic_vector(984,14),
		conv_std_logic_vector(990,14),
		conv_std_logic_vector(996,14),
		conv_std_logic_vector(1002,14),
		conv_std_logic_vector(1009,14),
		conv_std_logic_vector(1015,14),
		conv_std_logic_vector(1021,14),
		conv_std_logic_vector(1027,14),
		conv_std_logic_vector(1033,14),
		conv_std_logic_vector(1040,14),
		conv_std_logic_vector(1046,14),
		conv_std_logic_vector(1052,14),
		conv_std_logic_vector(1058,14),
		conv_std_logic_vector(1065,14),
		conv_std_logic_vector(1071,14),
		conv_std_logic_vector(1077,14),
		conv_std_logic_vector(1083,14),
		conv_std_logic_vector(1090,14),
		conv_std_logic_vector(1096,14),
		conv_std_logic_vector(1102,14),
		conv_std_logic_vector(1108,14),
		conv_std_logic_vector(1114,14),
		conv_std_logic_vector(1121,14),
		conv_std_logic_vector(1127,14),
		conv_std_logic_vector(1133,14),
		conv_std_logic_vector(1139,14),
		conv_std_logic_vector(1146,14),
		conv_std_logic_vector(1152,14),
		conv_std_logic_vector(1158,14),
		conv_std_logic_vector(1164,14),
		conv_std_logic_vector(1170,14),
		conv_std_logic_vector(1177,14),
		conv_std_logic_vector(1183,14),
		conv_std_logic_vector(1189,14),
		conv_std_logic_vector(1195,14),
		conv_std_logic_vector(1202,14),
		conv_std_logic_vector(1208,14),
		conv_std_logic_vector(1214,14),
		conv_std_logic_vector(1220,14),
		conv_std_logic_vector(1226,14),
		conv_std_logic_vector(1233,14),
		conv_std_logic_vector(1239,14),
		conv_std_logic_vector(1245,14),
		conv_std_logic_vector(1251,14),
		conv_std_logic_vector(1257,14),
		conv_std_logic_vector(1264,14),
		conv_std_logic_vector(1270,14),
		conv_std_logic_vector(1276,14),
		conv_std_logic_vector(1282,14),
		conv_std_logic_vector(1288,14),
		conv_std_logic_vector(1295,14),
		conv_std_logic_vector(1301,14),
		conv_std_logic_vector(1307,14),
		conv_std_logic_vector(1313,14),
		conv_std_logic_vector(1319,14),
		conv_std_logic_vector(1326,14),
		conv_std_logic_vector(1332,14),
		conv_std_logic_vector(1338,14),
		conv_std_logic_vector(1344,14),
		conv_std_logic_vector(1350,14),
		conv_std_logic_vector(1357,14),
		conv_std_logic_vector(1363,14),
		conv_std_logic_vector(1369,14),
		conv_std_logic_vector(1375,14),
		conv_std_logic_vector(1381,14),
		conv_std_logic_vector(1388,14),
		conv_std_logic_vector(1394,14),
		conv_std_logic_vector(1400,14),
		conv_std_logic_vector(1406,14),
		conv_std_logic_vector(1412,14),
		conv_std_logic_vector(1419,14),
		conv_std_logic_vector(1425,14),
		conv_std_logic_vector(1431,14),
		conv_std_logic_vector(1437,14),
		conv_std_logic_vector(1443,14),
		conv_std_logic_vector(1450,14),
		conv_std_logic_vector(1456,14),
		conv_std_logic_vector(1462,14),
		conv_std_logic_vector(1468,14),
		conv_std_logic_vector(1474,14),
		conv_std_logic_vector(1480,14),
		conv_std_logic_vector(1487,14),
		conv_std_logic_vector(1493,14),
		conv_std_logic_vector(1499,14),
		conv_std_logic_vector(1505,14),
		conv_std_logic_vector(1511,14),
		conv_std_logic_vector(1517,14),
		conv_std_logic_vector(1524,14),
		conv_std_logic_vector(1530,14),
		conv_std_logic_vector(1536,14),
		conv_std_logic_vector(1542,14),
		conv_std_logic_vector(1548,14),
		conv_std_logic_vector(1555,14),
		conv_std_logic_vector(1561,14),
		conv_std_logic_vector(1567,14),
		conv_std_logic_vector(1573,14),
		conv_std_logic_vector(1579,14),
		conv_std_logic_vector(1585,14),
		conv_std_logic_vector(1592,14),
		conv_std_logic_vector(1598,14),
		conv_std_logic_vector(1604,14),
		conv_std_logic_vector(1610,14),
		conv_std_logic_vector(1616,14),
		conv_std_logic_vector(1622,14),
		conv_std_logic_vector(1628,14),
		conv_std_logic_vector(1635,14),
		conv_std_logic_vector(1641,14),
		conv_std_logic_vector(1647,14),
		conv_std_logic_vector(1653,14),
		conv_std_logic_vector(1659,14),
		conv_std_logic_vector(1665,14),
		conv_std_logic_vector(1672,14),
		conv_std_logic_vector(1678,14),
		conv_std_logic_vector(1684,14),
		conv_std_logic_vector(1690,14),
		conv_std_logic_vector(1696,14),
		conv_std_logic_vector(1702,14),
		conv_std_logic_vector(1708,14),
		conv_std_logic_vector(1715,14),
		conv_std_logic_vector(1721,14),
		conv_std_logic_vector(1727,14),
		conv_std_logic_vector(1733,14),
		conv_std_logic_vector(1739,14),
		conv_std_logic_vector(1745,14),
		conv_std_logic_vector(1751,14),
		conv_std_logic_vector(1758,14),
		conv_std_logic_vector(1764,14),
		conv_std_logic_vector(1770,14),
		conv_std_logic_vector(1776,14),
		conv_std_logic_vector(1782,14),
		conv_std_logic_vector(1788,14),
		conv_std_logic_vector(1794,14),
		conv_std_logic_vector(1801,14),
		conv_std_logic_vector(1807,14),
		conv_std_logic_vector(1813,14),
		conv_std_logic_vector(1819,14),
		conv_std_logic_vector(1825,14),
		conv_std_logic_vector(1831,14),
		conv_std_logic_vector(1837,14),
		conv_std_logic_vector(1843,14),
		conv_std_logic_vector(1850,14),
		conv_std_logic_vector(1856,14),
		conv_std_logic_vector(1862,14),
		conv_std_logic_vector(1868,14),
		conv_std_logic_vector(1874,14),
		conv_std_logic_vector(1880,14),
		conv_std_logic_vector(1886,14),
		conv_std_logic_vector(1892,14),
		conv_std_logic_vector(1898,14),
		conv_std_logic_vector(1905,14),
		conv_std_logic_vector(1911,14),
		conv_std_logic_vector(1917,14),
		conv_std_logic_vector(1923,14),
		conv_std_logic_vector(1929,14),
		conv_std_logic_vector(1935,14),
		conv_std_logic_vector(1941,14),
		conv_std_logic_vector(1947,14),
		conv_std_logic_vector(1953,14),
		conv_std_logic_vector(1960,14),
		conv_std_logic_vector(1966,14),
		conv_std_logic_vector(1972,14),
		conv_std_logic_vector(1978,14),
		conv_std_logic_vector(1984,14),
		conv_std_logic_vector(1990,14),
		conv_std_logic_vector(1996,14),
		conv_std_logic_vector(2002,14),
		conv_std_logic_vector(2008,14),
		conv_std_logic_vector(2014,14),
		conv_std_logic_vector(2020,14),
		conv_std_logic_vector(2027,14),
		conv_std_logic_vector(2033,14),
		conv_std_logic_vector(2039,14),
		conv_std_logic_vector(2045,14),
		conv_std_logic_vector(2051,14),
		conv_std_logic_vector(2057,14),
		conv_std_logic_vector(2063,14),
		conv_std_logic_vector(2069,14),
		conv_std_logic_vector(2075,14),
		conv_std_logic_vector(2081,14),
		conv_std_logic_vector(2087,14),
		conv_std_logic_vector(2093,14),
		conv_std_logic_vector(2100,14),
		conv_std_logic_vector(2106,14),
		conv_std_logic_vector(2112,14),
		conv_std_logic_vector(2118,14),
		conv_std_logic_vector(2124,14),
		conv_std_logic_vector(2130,14),
		conv_std_logic_vector(2136,14),
		conv_std_logic_vector(2142,14),
		conv_std_logic_vector(2148,14),
		conv_std_logic_vector(2154,14),
		conv_std_logic_vector(2160,14),
		conv_std_logic_vector(2166,14),
		conv_std_logic_vector(2172,14),
		conv_std_logic_vector(2178,14),
		conv_std_logic_vector(2184,14),
		conv_std_logic_vector(2190,14),
		conv_std_logic_vector(2197,14),
		conv_std_logic_vector(2203,14),
		conv_std_logic_vector(2209,14),
		conv_std_logic_vector(2215,14),
		conv_std_logic_vector(2221,14),
		conv_std_logic_vector(2227,14),
		conv_std_logic_vector(2233,14),
		conv_std_logic_vector(2239,14),
		conv_std_logic_vector(2245,14),
		conv_std_logic_vector(2251,14),
		conv_std_logic_vector(2257,14),
		conv_std_logic_vector(2263,14),
		conv_std_logic_vector(2269,14),
		conv_std_logic_vector(2275,14),
		conv_std_logic_vector(2281,14),
		conv_std_logic_vector(2287,14),
		conv_std_logic_vector(2293,14),
		conv_std_logic_vector(2299,14),
		conv_std_logic_vector(2305,14),
		conv_std_logic_vector(2311,14),
		conv_std_logic_vector(2317,14),
		conv_std_logic_vector(2323,14),
		conv_std_logic_vector(2329,14),
		conv_std_logic_vector(2335,14),
		conv_std_logic_vector(2341,14),
		conv_std_logic_vector(2347,14),
		conv_std_logic_vector(2353,14),
		conv_std_logic_vector(2359,14),
		conv_std_logic_vector(2365,14),
		conv_std_logic_vector(2371,14),
		conv_std_logic_vector(2378,14),
		conv_std_logic_vector(2384,14),
		conv_std_logic_vector(2390,14),
		conv_std_logic_vector(2396,14),
		conv_std_logic_vector(2402,14),
		conv_std_logic_vector(2408,14),
		conv_std_logic_vector(2414,14),
		conv_std_logic_vector(2420,14),
		conv_std_logic_vector(2426,14),
		conv_std_logic_vector(2432,14),
		conv_std_logic_vector(2438,14),
		conv_std_logic_vector(2444,14),
		conv_std_logic_vector(2450,14),
		conv_std_logic_vector(2456,14),
		conv_std_logic_vector(2462,14),
		conv_std_logic_vector(2468,14),
		conv_std_logic_vector(2474,14),
		conv_std_logic_vector(2480,14),
		conv_std_logic_vector(2486,14),
		conv_std_logic_vector(2491,14),
		conv_std_logic_vector(2497,14),
		conv_std_logic_vector(2503,14),
		conv_std_logic_vector(2509,14),
		conv_std_logic_vector(2515,14),
		conv_std_logic_vector(2521,14),
		conv_std_logic_vector(2527,14),
		conv_std_logic_vector(2533,14),
		conv_std_logic_vector(2539,14),
		conv_std_logic_vector(2545,14),
		conv_std_logic_vector(2551,14),
		conv_std_logic_vector(2557,14),
		conv_std_logic_vector(2563,14),
		conv_std_logic_vector(2569,14),
		conv_std_logic_vector(2575,14),
		conv_std_logic_vector(2581,14),
		conv_std_logic_vector(2587,14),
		conv_std_logic_vector(2593,14),
		conv_std_logic_vector(2599,14),
		conv_std_logic_vector(2605,14),
		conv_std_logic_vector(2611,14),
		conv_std_logic_vector(2617,14),
		conv_std_logic_vector(2623,14),
		conv_std_logic_vector(2629,14),
		conv_std_logic_vector(2635,14),
		conv_std_logic_vector(2641,14),
		conv_std_logic_vector(2647,14),
		conv_std_logic_vector(2653,14),
		conv_std_logic_vector(2658,14),
		conv_std_logic_vector(2664,14),
		conv_std_logic_vector(2670,14),
		conv_std_logic_vector(2676,14),
		conv_std_logic_vector(2682,14),
		conv_std_logic_vector(2688,14),
		conv_std_logic_vector(2694,14),
		conv_std_logic_vector(2700,14),
		conv_std_logic_vector(2706,14),
		conv_std_logic_vector(2712,14),
		conv_std_logic_vector(2718,14),
		conv_std_logic_vector(2724,14),
		conv_std_logic_vector(2730,14),
		conv_std_logic_vector(2736,14),
		conv_std_logic_vector(2742,14),
		conv_std_logic_vector(2747,14),
		conv_std_logic_vector(2753,14),
		conv_std_logic_vector(2759,14),
		conv_std_logic_vector(2765,14),
		conv_std_logic_vector(2771,14),
		conv_std_logic_vector(2777,14),
		conv_std_logic_vector(2783,14),
		conv_std_logic_vector(2789,14),
		conv_std_logic_vector(2795,14),
		conv_std_logic_vector(2801,14),
		conv_std_logic_vector(2807,14),
		conv_std_logic_vector(2812,14),
		conv_std_logic_vector(2818,14),
		conv_std_logic_vector(2824,14),
		conv_std_logic_vector(2830,14),
		conv_std_logic_vector(2836,14),
		conv_std_logic_vector(2842,14),
		conv_std_logic_vector(2848,14),
		conv_std_logic_vector(2854,14),
		conv_std_logic_vector(2860,14),
		conv_std_logic_vector(2866,14),
		conv_std_logic_vector(2871,14),
		conv_std_logic_vector(2877,14),
		conv_std_logic_vector(2883,14),
		conv_std_logic_vector(2889,14),
		conv_std_logic_vector(2895,14),
		conv_std_logic_vector(2901,14),
		conv_std_logic_vector(2907,14),
		conv_std_logic_vector(2913,14),
		conv_std_logic_vector(2918,14),
		conv_std_logic_vector(2924,14),
		conv_std_logic_vector(2930,14),
		conv_std_logic_vector(2936,14),
		conv_std_logic_vector(2942,14),
		conv_std_logic_vector(2948,14),
		conv_std_logic_vector(2954,14),
		conv_std_logic_vector(2959,14),
		conv_std_logic_vector(2965,14),
		conv_std_logic_vector(2971,14),
		conv_std_logic_vector(2977,14),
		conv_std_logic_vector(2983,14),
		conv_std_logic_vector(2989,14),
		conv_std_logic_vector(2995,14),
		conv_std_logic_vector(3000,14),
		conv_std_logic_vector(3006,14),
		conv_std_logic_vector(3012,14),
		conv_std_logic_vector(3018,14),
		conv_std_logic_vector(3024,14),
		conv_std_logic_vector(3030,14),
		conv_std_logic_vector(3035,14),
		conv_std_logic_vector(3041,14),
		conv_std_logic_vector(3047,14),
		conv_std_logic_vector(3053,14),
		conv_std_logic_vector(3059,14),
		conv_std_logic_vector(3065,14),
		conv_std_logic_vector(3070,14),
		conv_std_logic_vector(3076,14),
		conv_std_logic_vector(3082,14),
		conv_std_logic_vector(3088,14),
		conv_std_logic_vector(3094,14),
		conv_std_logic_vector(3100,14),
		conv_std_logic_vector(3105,14),
		conv_std_logic_vector(3111,14),
		conv_std_logic_vector(3117,14),
		conv_std_logic_vector(3123,14),
		conv_std_logic_vector(3129,14),
		conv_std_logic_vector(3134,14),
		conv_std_logic_vector(3140,14),
		conv_std_logic_vector(3146,14),
		conv_std_logic_vector(3152,14),
		conv_std_logic_vector(3158,14),
		conv_std_logic_vector(3163,14),
		conv_std_logic_vector(3169,14),
		conv_std_logic_vector(3175,14),
		conv_std_logic_vector(3181,14),
		conv_std_logic_vector(3187,14),
		conv_std_logic_vector(3192,14),
		conv_std_logic_vector(3198,14),
		conv_std_logic_vector(3204,14),
		conv_std_logic_vector(3210,14),
		conv_std_logic_vector(3216,14),
		conv_std_logic_vector(3221,14),
		conv_std_logic_vector(3227,14),
		conv_std_logic_vector(3233,14),
		conv_std_logic_vector(3239,14),
		conv_std_logic_vector(3244,14),
		conv_std_logic_vector(3250,14),
		conv_std_logic_vector(3256,14),
		conv_std_logic_vector(3262,14),
		conv_std_logic_vector(3267,14),
		conv_std_logic_vector(3273,14),
		conv_std_logic_vector(3279,14),
		conv_std_logic_vector(3285,14),
		conv_std_logic_vector(3290,14),
		conv_std_logic_vector(3296,14),
		conv_std_logic_vector(3302,14),
		conv_std_logic_vector(3308,14),
		conv_std_logic_vector(3313,14),
		conv_std_logic_vector(3319,14),
		conv_std_logic_vector(3325,14),
		conv_std_logic_vector(3331,14),
		conv_std_logic_vector(3336,14),
		conv_std_logic_vector(3342,14),
		conv_std_logic_vector(3348,14),
		conv_std_logic_vector(3354,14),
		conv_std_logic_vector(3359,14),
		conv_std_logic_vector(3365,14),
		conv_std_logic_vector(3371,14),
		conv_std_logic_vector(3377,14),
		conv_std_logic_vector(3382,14),
		conv_std_logic_vector(3388,14),
		conv_std_logic_vector(3394,14),
		conv_std_logic_vector(3399,14),
		conv_std_logic_vector(3405,14),
		conv_std_logic_vector(3411,14),
		conv_std_logic_vector(3417,14),
		conv_std_logic_vector(3422,14),
		conv_std_logic_vector(3428,14),
		conv_std_logic_vector(3434,14),
		conv_std_logic_vector(3439,14),
		conv_std_logic_vector(3445,14),
		conv_std_logic_vector(3451,14),
		conv_std_logic_vector(3457,14),
		conv_std_logic_vector(3462,14),
		conv_std_logic_vector(3468,14),
		conv_std_logic_vector(3474,14),
		conv_std_logic_vector(3479,14),
		conv_std_logic_vector(3485,14),
		conv_std_logic_vector(3491,14),
		conv_std_logic_vector(3496,14),
		conv_std_logic_vector(3502,14),
		conv_std_logic_vector(3508,14),
		conv_std_logic_vector(3513,14),
		conv_std_logic_vector(3519,14),
		conv_std_logic_vector(3525,14),
		conv_std_logic_vector(3530,14),
		conv_std_logic_vector(3536,14),
		conv_std_logic_vector(3542,14),
		conv_std_logic_vector(3547,14),
		conv_std_logic_vector(3553,14),
		conv_std_logic_vector(3559,14),
		conv_std_logic_vector(3564,14),
		conv_std_logic_vector(3570,14),
		conv_std_logic_vector(3576,14),
		conv_std_logic_vector(3581,14),
		conv_std_logic_vector(3587,14),
		conv_std_logic_vector(3593,14),
		conv_std_logic_vector(3598,14),
		conv_std_logic_vector(3604,14),
		conv_std_logic_vector(3610,14),
		conv_std_logic_vector(3615,14),
		conv_std_logic_vector(3621,14),
		conv_std_logic_vector(3626,14),
		conv_std_logic_vector(3632,14),
		conv_std_logic_vector(3638,14),
		conv_std_logic_vector(3643,14),
		conv_std_logic_vector(3649,14),
		conv_std_logic_vector(3655,14),
		conv_std_logic_vector(3660,14),
		conv_std_logic_vector(3666,14),
		conv_std_logic_vector(3671,14),
		conv_std_logic_vector(3677,14),
		conv_std_logic_vector(3683,14),
		conv_std_logic_vector(3688,14),
		conv_std_logic_vector(3694,14),
		conv_std_logic_vector(3700,14),
		conv_std_logic_vector(3705,14),
		conv_std_logic_vector(3711,14),
		conv_std_logic_vector(3716,14),
		conv_std_logic_vector(3722,14),
		conv_std_logic_vector(3728,14),
		conv_std_logic_vector(3733,14),
		conv_std_logic_vector(3739,14),
		conv_std_logic_vector(3744,14),
		conv_std_logic_vector(3750,14),
		conv_std_logic_vector(3755,14),
		conv_std_logic_vector(3761,14),
		conv_std_logic_vector(3767,14),
		conv_std_logic_vector(3772,14),
		conv_std_logic_vector(3778,14),
		conv_std_logic_vector(3783,14),
		conv_std_logic_vector(3789,14),
		conv_std_logic_vector(3795,14),
		conv_std_logic_vector(3800,14),
		conv_std_logic_vector(3806,14),
		conv_std_logic_vector(3811,14),
		conv_std_logic_vector(3817,14),
		conv_std_logic_vector(3822,14),
		conv_std_logic_vector(3828,14),
		conv_std_logic_vector(3833,14),
		conv_std_logic_vector(3839,14),
		conv_std_logic_vector(3845,14),
		conv_std_logic_vector(3850,14),
		conv_std_logic_vector(3856,14),
		conv_std_logic_vector(3861,14),
		conv_std_logic_vector(3867,14),
		conv_std_logic_vector(3872,14),
		conv_std_logic_vector(3878,14),
		conv_std_logic_vector(3883,14),
		conv_std_logic_vector(3889,14),
		conv_std_logic_vector(3894,14),
		conv_std_logic_vector(3900,14),
		conv_std_logic_vector(3905,14),
		conv_std_logic_vector(3911,14),
		conv_std_logic_vector(3916,14),
		conv_std_logic_vector(3922,14),
		conv_std_logic_vector(3928,14),
		conv_std_logic_vector(3933,14),
		conv_std_logic_vector(3939,14),
		conv_std_logic_vector(3944,14),
		conv_std_logic_vector(3950,14),
		conv_std_logic_vector(3955,14),
		conv_std_logic_vector(3961,14),
		conv_std_logic_vector(3966,14),
		conv_std_logic_vector(3972,14),
		conv_std_logic_vector(3977,14),
		conv_std_logic_vector(3983,14),
		conv_std_logic_vector(3988,14),
		conv_std_logic_vector(3994,14),
		conv_std_logic_vector(3999,14),
		conv_std_logic_vector(4004,14),
		conv_std_logic_vector(4010,14),
		conv_std_logic_vector(4015,14),
		conv_std_logic_vector(4021,14),
		conv_std_logic_vector(4026,14),
		conv_std_logic_vector(4032,14),
		conv_std_logic_vector(4037,14),
		conv_std_logic_vector(4043,14),
		conv_std_logic_vector(4048,14),
		conv_std_logic_vector(4054,14),
		conv_std_logic_vector(4059,14),
		conv_std_logic_vector(4065,14),
		conv_std_logic_vector(4070,14),
		conv_std_logic_vector(4076,14),
		conv_std_logic_vector(4081,14),
		conv_std_logic_vector(4086,14),
		conv_std_logic_vector(4092,14),
		conv_std_logic_vector(4097,14),
		conv_std_logic_vector(4103,14),
		conv_std_logic_vector(4108,14),
		conv_std_logic_vector(4114,14),
		conv_std_logic_vector(4119,14),
		conv_std_logic_vector(4124,14),
		conv_std_logic_vector(4130,14),
		conv_std_logic_vector(4135,14),
		conv_std_logic_vector(4141,14),
		conv_std_logic_vector(4146,14),
		conv_std_logic_vector(4152,14),
		conv_std_logic_vector(4157,14),
		conv_std_logic_vector(4162,14),
		conv_std_logic_vector(4168,14),
		conv_std_logic_vector(4173,14),
		conv_std_logic_vector(4179,14),
		conv_std_logic_vector(4184,14),
		conv_std_logic_vector(4189,14),
		conv_std_logic_vector(4195,14),
		conv_std_logic_vector(4200,14),
		conv_std_logic_vector(4206,14),
		conv_std_logic_vector(4211,14),
		conv_std_logic_vector(4216,14),
		conv_std_logic_vector(4222,14),
		conv_std_logic_vector(4227,14),
		conv_std_logic_vector(4233,14),
		conv_std_logic_vector(4238,14),
		conv_std_logic_vector(4243,14),
		conv_std_logic_vector(4249,14),
		conv_std_logic_vector(4254,14),
		conv_std_logic_vector(4259,14),
		conv_std_logic_vector(4265,14),
		conv_std_logic_vector(4270,14),
		conv_std_logic_vector(4276,14),
		conv_std_logic_vector(4281,14),
		conv_std_logic_vector(4286,14),
		conv_std_logic_vector(4292,14),
		conv_std_logic_vector(4297,14),
		conv_std_logic_vector(4302,14),
		conv_std_logic_vector(4308,14),
		conv_std_logic_vector(4313,14),
		conv_std_logic_vector(4318,14),
		conv_std_logic_vector(4324,14),
		conv_std_logic_vector(4329,14),
		conv_std_logic_vector(4334,14),
		conv_std_logic_vector(4340,14),
		conv_std_logic_vector(4345,14),
		conv_std_logic_vector(4350,14),
		conv_std_logic_vector(4356,14),
		conv_std_logic_vector(4361,14),
		conv_std_logic_vector(4366,14),
		conv_std_logic_vector(4372,14),
		conv_std_logic_vector(4377,14),
		conv_std_logic_vector(4382,14),
		conv_std_logic_vector(4388,14),
		conv_std_logic_vector(4393,14),
		conv_std_logic_vector(4398,14),
		conv_std_logic_vector(4403,14),
		conv_std_logic_vector(4409,14),
		conv_std_logic_vector(4414,14),
		conv_std_logic_vector(4419,14),
		conv_std_logic_vector(4425,14),
		conv_std_logic_vector(4430,14),
		conv_std_logic_vector(4435,14),
		conv_std_logic_vector(4440,14),
		conv_std_logic_vector(4446,14),
		conv_std_logic_vector(4451,14),
		conv_std_logic_vector(4456,14),
		conv_std_logic_vector(4462,14),
		conv_std_logic_vector(4467,14),
		conv_std_logic_vector(4472,14),
		conv_std_logic_vector(4477,14),
		conv_std_logic_vector(4483,14),
		conv_std_logic_vector(4488,14),
		conv_std_logic_vector(4493,14),
		conv_std_logic_vector(4498,14),
		conv_std_logic_vector(4504,14),
		conv_std_logic_vector(4509,14),
		conv_std_logic_vector(4514,14),
		conv_std_logic_vector(4519,14),
		conv_std_logic_vector(4525,14),
		conv_std_logic_vector(4530,14),
		conv_std_logic_vector(4535,14),
		conv_std_logic_vector(4540,14),
		conv_std_logic_vector(4546,14),
		conv_std_logic_vector(4551,14),
		conv_std_logic_vector(4556,14),
		conv_std_logic_vector(4561,14),
		conv_std_logic_vector(4566,14),
		conv_std_logic_vector(4572,14),
		conv_std_logic_vector(4577,14),
		conv_std_logic_vector(4582,14),
		conv_std_logic_vector(4587,14),
		conv_std_logic_vector(4592,14),
		conv_std_logic_vector(4598,14),
		conv_std_logic_vector(4603,14),
		conv_std_logic_vector(4608,14),
		conv_std_logic_vector(4613,14),
		conv_std_logic_vector(4618,14),
		conv_std_logic_vector(4624,14),
		conv_std_logic_vector(4629,14),
		conv_std_logic_vector(4634,14),
		conv_std_logic_vector(4639,14),
		conv_std_logic_vector(4644,14),
		conv_std_logic_vector(4650,14),
		conv_std_logic_vector(4655,14),
		conv_std_logic_vector(4660,14),
		conv_std_logic_vector(4665,14),
		conv_std_logic_vector(4670,14),
		conv_std_logic_vector(4675,14),
		conv_std_logic_vector(4680,14),
		conv_std_logic_vector(4686,14),
		conv_std_logic_vector(4691,14),
		conv_std_logic_vector(4696,14),
		conv_std_logic_vector(4701,14),
		conv_std_logic_vector(4706,14),
		conv_std_logic_vector(4711,14),
		conv_std_logic_vector(4717,14),
		conv_std_logic_vector(4722,14),
		conv_std_logic_vector(4727,14),
		conv_std_logic_vector(4732,14),
		conv_std_logic_vector(4737,14),
		conv_std_logic_vector(4742,14),
		conv_std_logic_vector(4747,14),
		conv_std_logic_vector(4752,14),
		conv_std_logic_vector(4758,14),
		conv_std_logic_vector(4763,14),
		conv_std_logic_vector(4768,14),
		conv_std_logic_vector(4773,14),
		conv_std_logic_vector(4778,14),
		conv_std_logic_vector(4783,14),
		conv_std_logic_vector(4788,14),
		conv_std_logic_vector(4793,14),
		conv_std_logic_vector(4798,14),
		conv_std_logic_vector(4803,14),
		conv_std_logic_vector(4809,14),
		conv_std_logic_vector(4814,14),
		conv_std_logic_vector(4819,14),
		conv_std_logic_vector(4824,14),
		conv_std_logic_vector(4829,14),
		conv_std_logic_vector(4834,14),
		conv_std_logic_vector(4839,14),
		conv_std_logic_vector(4844,14),
		conv_std_logic_vector(4849,14),
		conv_std_logic_vector(4854,14),
		conv_std_logic_vector(4859,14),
		conv_std_logic_vector(4864,14),
		conv_std_logic_vector(4869,14),
		conv_std_logic_vector(4874,14),
		conv_std_logic_vector(4879,14),
		conv_std_logic_vector(4885,14),
		conv_std_logic_vector(4890,14),
		conv_std_logic_vector(4895,14),
		conv_std_logic_vector(4900,14),
		conv_std_logic_vector(4905,14),
		conv_std_logic_vector(4910,14),
		conv_std_logic_vector(4915,14),
		conv_std_logic_vector(4920,14),
		conv_std_logic_vector(4925,14),
		conv_std_logic_vector(4930,14),
		conv_std_logic_vector(4935,14),
		conv_std_logic_vector(4940,14),
		conv_std_logic_vector(4945,14),
		conv_std_logic_vector(4950,14),
		conv_std_logic_vector(4955,14),
		conv_std_logic_vector(4960,14),
		conv_std_logic_vector(4965,14),
		conv_std_logic_vector(4970,14),
		conv_std_logic_vector(4975,14),
		conv_std_logic_vector(4980,14),
		conv_std_logic_vector(4985,14),
		conv_std_logic_vector(4990,14),
		conv_std_logic_vector(4995,14),
		conv_std_logic_vector(5000,14),
		conv_std_logic_vector(5005,14),
		conv_std_logic_vector(5010,14),
		conv_std_logic_vector(5015,14),
		conv_std_logic_vector(5020,14),
		conv_std_logic_vector(5025,14),
		conv_std_logic_vector(5030,14),
		conv_std_logic_vector(5035,14),
		conv_std_logic_vector(5039,14),
		conv_std_logic_vector(5044,14),
		conv_std_logic_vector(5049,14),
		conv_std_logic_vector(5054,14),
		conv_std_logic_vector(5059,14),
		conv_std_logic_vector(5064,14),
		conv_std_logic_vector(5069,14),
		conv_std_logic_vector(5074,14),
		conv_std_logic_vector(5079,14),
		conv_std_logic_vector(5084,14),
		conv_std_logic_vector(5089,14),
		conv_std_logic_vector(5094,14),
		conv_std_logic_vector(5099,14),
		conv_std_logic_vector(5104,14),
		conv_std_logic_vector(5109,14),
		conv_std_logic_vector(5113,14),
		conv_std_logic_vector(5118,14),
		conv_std_logic_vector(5123,14),
		conv_std_logic_vector(5128,14),
		conv_std_logic_vector(5133,14),
		conv_std_logic_vector(5138,14),
		conv_std_logic_vector(5143,14),
		conv_std_logic_vector(5148,14),
		conv_std_logic_vector(5153,14),
		conv_std_logic_vector(5157,14),
		conv_std_logic_vector(5162,14),
		conv_std_logic_vector(5167,14),
		conv_std_logic_vector(5172,14),
		conv_std_logic_vector(5177,14),
		conv_std_logic_vector(5182,14),
		conv_std_logic_vector(5187,14),
		conv_std_logic_vector(5192,14),
		conv_std_logic_vector(5196,14),
		conv_std_logic_vector(5201,14),
		conv_std_logic_vector(5206,14),
		conv_std_logic_vector(5211,14),
		conv_std_logic_vector(5216,14),
		conv_std_logic_vector(5221,14),
		conv_std_logic_vector(5226,14),
		conv_std_logic_vector(5230,14),
		conv_std_logic_vector(5235,14),
		conv_std_logic_vector(5240,14),
		conv_std_logic_vector(5245,14),
		conv_std_logic_vector(5250,14),
		conv_std_logic_vector(5255,14),
		conv_std_logic_vector(5259,14),
		conv_std_logic_vector(5264,14),
		conv_std_logic_vector(5269,14),
		conv_std_logic_vector(5274,14),
		conv_std_logic_vector(5279,14),
		conv_std_logic_vector(5283,14),
		conv_std_logic_vector(5288,14),
		conv_std_logic_vector(5293,14),
		conv_std_logic_vector(5298,14),
		conv_std_logic_vector(5303,14),
		conv_std_logic_vector(5307,14),
		conv_std_logic_vector(5312,14),
		conv_std_logic_vector(5317,14),
		conv_std_logic_vector(5322,14),
		conv_std_logic_vector(5326,14),
		conv_std_logic_vector(5331,14),
		conv_std_logic_vector(5336,14),
		conv_std_logic_vector(5341,14),
		conv_std_logic_vector(5346,14),
		conv_std_logic_vector(5350,14),
		conv_std_logic_vector(5355,14),
		conv_std_logic_vector(5360,14),
		conv_std_logic_vector(5365,14),
		conv_std_logic_vector(5369,14),
		conv_std_logic_vector(5374,14),
		conv_std_logic_vector(5379,14),
		conv_std_logic_vector(5384,14),
		conv_std_logic_vector(5388,14),
		conv_std_logic_vector(5393,14),
		conv_std_logic_vector(5398,14),
		conv_std_logic_vector(5402,14),
		conv_std_logic_vector(5407,14),
		conv_std_logic_vector(5412,14),
		conv_std_logic_vector(5417,14),
		conv_std_logic_vector(5421,14),
		conv_std_logic_vector(5426,14),
		conv_std_logic_vector(5431,14),
		conv_std_logic_vector(5435,14),
		conv_std_logic_vector(5440,14),
		conv_std_logic_vector(5445,14),
		conv_std_logic_vector(5450,14),
		conv_std_logic_vector(5454,14),
		conv_std_logic_vector(5459,14),
		conv_std_logic_vector(5464,14),
		conv_std_logic_vector(5468,14),
		conv_std_logic_vector(5473,14),
		conv_std_logic_vector(5478,14),
		conv_std_logic_vector(5482,14),
		conv_std_logic_vector(5487,14),
		conv_std_logic_vector(5492,14),
		conv_std_logic_vector(5496,14),
		conv_std_logic_vector(5501,14),
		conv_std_logic_vector(5506,14),
		conv_std_logic_vector(5510,14),
		conv_std_logic_vector(5515,14),
		conv_std_logic_vector(5520,14),
		conv_std_logic_vector(5524,14),
		conv_std_logic_vector(5529,14),
		conv_std_logic_vector(5533,14),
		conv_std_logic_vector(5538,14),
		conv_std_logic_vector(5543,14),
		conv_std_logic_vector(5547,14),
		conv_std_logic_vector(5552,14),
		conv_std_logic_vector(5557,14),
		conv_std_logic_vector(5561,14),
		conv_std_logic_vector(5566,14),
		conv_std_logic_vector(5570,14),
		conv_std_logic_vector(5575,14),
		conv_std_logic_vector(5580,14),
		conv_std_logic_vector(5584,14),
		conv_std_logic_vector(5589,14),
		conv_std_logic_vector(5593,14),
		conv_std_logic_vector(5598,14),
		conv_std_logic_vector(5603,14),
		conv_std_logic_vector(5607,14),
		conv_std_logic_vector(5612,14),
		conv_std_logic_vector(5616,14),
		conv_std_logic_vector(5621,14),
		conv_std_logic_vector(5625,14),
		conv_std_logic_vector(5630,14),
		conv_std_logic_vector(5635,14),
		conv_std_logic_vector(5639,14),
		conv_std_logic_vector(5644,14),
		conv_std_logic_vector(5648,14),
		conv_std_logic_vector(5653,14),
		conv_std_logic_vector(5657,14),
		conv_std_logic_vector(5662,14),
		conv_std_logic_vector(5666,14),
		conv_std_logic_vector(5671,14),
		conv_std_logic_vector(5675,14),
		conv_std_logic_vector(5680,14),
		conv_std_logic_vector(5685,14),
		conv_std_logic_vector(5689,14),
		conv_std_logic_vector(5694,14),
		conv_std_logic_vector(5698,14),
		conv_std_logic_vector(5703,14),
		conv_std_logic_vector(5707,14),
		conv_std_logic_vector(5712,14),
		conv_std_logic_vector(5716,14),
		conv_std_logic_vector(5721,14),
		conv_std_logic_vector(5725,14),
		conv_std_logic_vector(5730,14),
		conv_std_logic_vector(5734,14),
		conv_std_logic_vector(5739,14),
		conv_std_logic_vector(5743,14),
		conv_std_logic_vector(5748,14),
		conv_std_logic_vector(5752,14),
		conv_std_logic_vector(5756,14),
		conv_std_logic_vector(5761,14),
		conv_std_logic_vector(5765,14),
		conv_std_logic_vector(5770,14),
		conv_std_logic_vector(5774,14),
		conv_std_logic_vector(5779,14),
		conv_std_logic_vector(5783,14),
		conv_std_logic_vector(5788,14),
		conv_std_logic_vector(5792,14),
		conv_std_logic_vector(5797,14),
		conv_std_logic_vector(5801,14),
		conv_std_logic_vector(5805,14),
		conv_std_logic_vector(5810,14),
		conv_std_logic_vector(5814,14),
		conv_std_logic_vector(5819,14),
		conv_std_logic_vector(5823,14),
		conv_std_logic_vector(5828,14),
		conv_std_logic_vector(5832,14),
		conv_std_logic_vector(5836,14),
		conv_std_logic_vector(5841,14),
		conv_std_logic_vector(5845,14),
		conv_std_logic_vector(5850,14),
		conv_std_logic_vector(5854,14),
		conv_std_logic_vector(5858,14),
		conv_std_logic_vector(5863,14),
		conv_std_logic_vector(5867,14),
		conv_std_logic_vector(5872,14),
		conv_std_logic_vector(5876,14),
		conv_std_logic_vector(5880,14),
		conv_std_logic_vector(5885,14),
		conv_std_logic_vector(5889,14),
		conv_std_logic_vector(5893,14),
		conv_std_logic_vector(5898,14),
		conv_std_logic_vector(5902,14),
		conv_std_logic_vector(5906,14),
		conv_std_logic_vector(5911,14),
		conv_std_logic_vector(5915,14),
		conv_std_logic_vector(5920,14),
		conv_std_logic_vector(5924,14),
		conv_std_logic_vector(5928,14),
		conv_std_logic_vector(5933,14),
		conv_std_logic_vector(5937,14),
		conv_std_logic_vector(5941,14),
		conv_std_logic_vector(5946,14),
		conv_std_logic_vector(5950,14),
		conv_std_logic_vector(5954,14),
		conv_std_logic_vector(5958,14),
		conv_std_logic_vector(5963,14),
		conv_std_logic_vector(5967,14),
		conv_std_logic_vector(5971,14),
		conv_std_logic_vector(5976,14),
		conv_std_logic_vector(5980,14),
		conv_std_logic_vector(5984,14),
		conv_std_logic_vector(5989,14),
		conv_std_logic_vector(5993,14),
		conv_std_logic_vector(5997,14),
		conv_std_logic_vector(6001,14),
		conv_std_logic_vector(6006,14),
		conv_std_logic_vector(6010,14),
		conv_std_logic_vector(6014,14),
		conv_std_logic_vector(6018,14),
		conv_std_logic_vector(6023,14),
		conv_std_logic_vector(6027,14),
		conv_std_logic_vector(6031,14),
		conv_std_logic_vector(6036,14),
		conv_std_logic_vector(6040,14),
		conv_std_logic_vector(6044,14),
		conv_std_logic_vector(6048,14),
		conv_std_logic_vector(6052,14),
		conv_std_logic_vector(6057,14),
		conv_std_logic_vector(6061,14),
		conv_std_logic_vector(6065,14),
		conv_std_logic_vector(6069,14),
		conv_std_logic_vector(6074,14),
		conv_std_logic_vector(6078,14),
		conv_std_logic_vector(6082,14),
		conv_std_logic_vector(6086,14),
		conv_std_logic_vector(6090,14),
		conv_std_logic_vector(6095,14),
		conv_std_logic_vector(6099,14),
		conv_std_logic_vector(6103,14),
		conv_std_logic_vector(6107,14),
		conv_std_logic_vector(6111,14),
		conv_std_logic_vector(6116,14),
		conv_std_logic_vector(6120,14),
		conv_std_logic_vector(6124,14),
		conv_std_logic_vector(6128,14),
		conv_std_logic_vector(6132,14),
		conv_std_logic_vector(6136,14),
		conv_std_logic_vector(6141,14),
		conv_std_logic_vector(6145,14),
		conv_std_logic_vector(6149,14),
		conv_std_logic_vector(6153,14),
		conv_std_logic_vector(6157,14),
		conv_std_logic_vector(6161,14),
		conv_std_logic_vector(6165,14),
		conv_std_logic_vector(6170,14),
		conv_std_logic_vector(6174,14),
		conv_std_logic_vector(6178,14),
		conv_std_logic_vector(6182,14),
		conv_std_logic_vector(6186,14),
		conv_std_logic_vector(6190,14),
		conv_std_logic_vector(6194,14),
		conv_std_logic_vector(6198,14),
		conv_std_logic_vector(6203,14),
		conv_std_logic_vector(6207,14),
		conv_std_logic_vector(6211,14),
		conv_std_logic_vector(6215,14),
		conv_std_logic_vector(6219,14),
		conv_std_logic_vector(6223,14),
		conv_std_logic_vector(6227,14),
		conv_std_logic_vector(6231,14),
		conv_std_logic_vector(6235,14),
		conv_std_logic_vector(6239,14),
		conv_std_logic_vector(6243,14),
		conv_std_logic_vector(6247,14),
		conv_std_logic_vector(6252,14),
		conv_std_logic_vector(6256,14),
		conv_std_logic_vector(6260,14),
		conv_std_logic_vector(6264,14),
		conv_std_logic_vector(6268,14),
		conv_std_logic_vector(6272,14),
		conv_std_logic_vector(6276,14),
		conv_std_logic_vector(6280,14),
		conv_std_logic_vector(6284,14),
		conv_std_logic_vector(6288,14),
		conv_std_logic_vector(6292,14),
		conv_std_logic_vector(6296,14),
		conv_std_logic_vector(6300,14),
		conv_std_logic_vector(6304,14),
		conv_std_logic_vector(6308,14),
		conv_std_logic_vector(6312,14),
		conv_std_logic_vector(6316,14),
		conv_std_logic_vector(6320,14),
		conv_std_logic_vector(6324,14),
		conv_std_logic_vector(6328,14),
		conv_std_logic_vector(6332,14),
		conv_std_logic_vector(6336,14),
		conv_std_logic_vector(6340,14),
		conv_std_logic_vector(6344,14),
		conv_std_logic_vector(6348,14),
		conv_std_logic_vector(6352,14),
		conv_std_logic_vector(6356,14),
		conv_std_logic_vector(6360,14),
		conv_std_logic_vector(6364,14),
		conv_std_logic_vector(6368,14),
		conv_std_logic_vector(6372,14),
		conv_std_logic_vector(6376,14),
		conv_std_logic_vector(6380,14),
		conv_std_logic_vector(6384,14),
		conv_std_logic_vector(6387,14),
		conv_std_logic_vector(6391,14),
		conv_std_logic_vector(6395,14),
		conv_std_logic_vector(6399,14),
		conv_std_logic_vector(6403,14),
		conv_std_logic_vector(6407,14),
		conv_std_logic_vector(6411,14),
		conv_std_logic_vector(6415,14),
		conv_std_logic_vector(6419,14),
		conv_std_logic_vector(6423,14),
		conv_std_logic_vector(6427,14),
		conv_std_logic_vector(6430,14),
		conv_std_logic_vector(6434,14),
		conv_std_logic_vector(6438,14),
		conv_std_logic_vector(6442,14),
		conv_std_logic_vector(6446,14),
		conv_std_logic_vector(6450,14),
		conv_std_logic_vector(6454,14),
		conv_std_logic_vector(6458,14),
		conv_std_logic_vector(6461,14),
		conv_std_logic_vector(6465,14),
		conv_std_logic_vector(6469,14),
		conv_std_logic_vector(6473,14),
		conv_std_logic_vector(6477,14),
		conv_std_logic_vector(6481,14),
		conv_std_logic_vector(6485,14),
		conv_std_logic_vector(6488,14),
		conv_std_logic_vector(6492,14),
		conv_std_logic_vector(6496,14),
		conv_std_logic_vector(6500,14),
		conv_std_logic_vector(6504,14),
		conv_std_logic_vector(6508,14),
		conv_std_logic_vector(6511,14),
		conv_std_logic_vector(6515,14),
		conv_std_logic_vector(6519,14),
		conv_std_logic_vector(6523,14),
		conv_std_logic_vector(6527,14),
		conv_std_logic_vector(6530,14),
		conv_std_logic_vector(6534,14),
		conv_std_logic_vector(6538,14),
		conv_std_logic_vector(6542,14),
		conv_std_logic_vector(6546,14),
		conv_std_logic_vector(6549,14),
		conv_std_logic_vector(6553,14),
		conv_std_logic_vector(6557,14),
		conv_std_logic_vector(6561,14),
		conv_std_logic_vector(6564,14),
		conv_std_logic_vector(6568,14),
		conv_std_logic_vector(6572,14),
		conv_std_logic_vector(6576,14),
		conv_std_logic_vector(6579,14),
		conv_std_logic_vector(6583,14),
		conv_std_logic_vector(6587,14),
		conv_std_logic_vector(6591,14),
		conv_std_logic_vector(6594,14),
		conv_std_logic_vector(6598,14),
		conv_std_logic_vector(6602,14),
		conv_std_logic_vector(6605,14),
		conv_std_logic_vector(6609,14),
		conv_std_logic_vector(6613,14),
		conv_std_logic_vector(6617,14),
		conv_std_logic_vector(6620,14),
		conv_std_logic_vector(6624,14),
		conv_std_logic_vector(6628,14),
		conv_std_logic_vector(6631,14),
		conv_std_logic_vector(6635,14),
		conv_std_logic_vector(6639,14),
		conv_std_logic_vector(6642,14),
		conv_std_logic_vector(6646,14),
		conv_std_logic_vector(6650,14),
		conv_std_logic_vector(6653,14),
		conv_std_logic_vector(6657,14),
		conv_std_logic_vector(6661,14),
		conv_std_logic_vector(6664,14),
		conv_std_logic_vector(6668,14),
		conv_std_logic_vector(6672,14),
		conv_std_logic_vector(6675,14),
		conv_std_logic_vector(6679,14),
		conv_std_logic_vector(6683,14),
		conv_std_logic_vector(6686,14),
		conv_std_logic_vector(6690,14),
		conv_std_logic_vector(6694,14),
		conv_std_logic_vector(6697,14),
		conv_std_logic_vector(6701,14),
		conv_std_logic_vector(6704,14),
		conv_std_logic_vector(6708,14),
		conv_std_logic_vector(6712,14),
		conv_std_logic_vector(6715,14),
		conv_std_logic_vector(6719,14),
		conv_std_logic_vector(6722,14),
		conv_std_logic_vector(6726,14),
		conv_std_logic_vector(6730,14),
		conv_std_logic_vector(6733,14),
		conv_std_logic_vector(6737,14),
		conv_std_logic_vector(6740,14),
		conv_std_logic_vector(6744,14),
		conv_std_logic_vector(6747,14),
		conv_std_logic_vector(6751,14),
		conv_std_logic_vector(6755,14),
		conv_std_logic_vector(6758,14),
		conv_std_logic_vector(6762,14),
		conv_std_logic_vector(6765,14),
		conv_std_logic_vector(6769,14),
		conv_std_logic_vector(6772,14),
		conv_std_logic_vector(6776,14),
		conv_std_logic_vector(6779,14),
		conv_std_logic_vector(6783,14),
		conv_std_logic_vector(6786,14),
		conv_std_logic_vector(6790,14),
		conv_std_logic_vector(6793,14),
		conv_std_logic_vector(6797,14),
		conv_std_logic_vector(6800,14),
		conv_std_logic_vector(6804,14),
		conv_std_logic_vector(6807,14),
		conv_std_logic_vector(6811,14),
		conv_std_logic_vector(6814,14),
		conv_std_logic_vector(6818,14),
		conv_std_logic_vector(6821,14),
		conv_std_logic_vector(6825,14),
		conv_std_logic_vector(6828,14),
		conv_std_logic_vector(6832,14),
		conv_std_logic_vector(6835,14),
		conv_std_logic_vector(6839,14),
		conv_std_logic_vector(6842,14),
		conv_std_logic_vector(6846,14),
		conv_std_logic_vector(6849,14),
		conv_std_logic_vector(6852,14),
		conv_std_logic_vector(6856,14),
		conv_std_logic_vector(6859,14),
		conv_std_logic_vector(6863,14),
		conv_std_logic_vector(6866,14),
		conv_std_logic_vector(6870,14),
		conv_std_logic_vector(6873,14),
		conv_std_logic_vector(6876,14),
		conv_std_logic_vector(6880,14),
		conv_std_logic_vector(6883,14),
		conv_std_logic_vector(6887,14),
		conv_std_logic_vector(6890,14),
		conv_std_logic_vector(6894,14),
		conv_std_logic_vector(6897,14),
		conv_std_logic_vector(6900,14),
		conv_std_logic_vector(6904,14),
		conv_std_logic_vector(6907,14),
		conv_std_logic_vector(6910,14),
		conv_std_logic_vector(6914,14),
		conv_std_logic_vector(6917,14),
		conv_std_logic_vector(6921,14),
		conv_std_logic_vector(6924,14),
		conv_std_logic_vector(6927,14),
		conv_std_logic_vector(6931,14),
		conv_std_logic_vector(6934,14),
		conv_std_logic_vector(6937,14),
		conv_std_logic_vector(6941,14),
		conv_std_logic_vector(6944,14),
		conv_std_logic_vector(6947,14),
		conv_std_logic_vector(6951,14),
		conv_std_logic_vector(6954,14),
		conv_std_logic_vector(6957,14),
		conv_std_logic_vector(6961,14),
		conv_std_logic_vector(6964,14),
		conv_std_logic_vector(6967,14),
		conv_std_logic_vector(6971,14),
		conv_std_logic_vector(6974,14),
		conv_std_logic_vector(6977,14),
		conv_std_logic_vector(6980,14),
		conv_std_logic_vector(6984,14),
		conv_std_logic_vector(6987,14),
		conv_std_logic_vector(6990,14),
		conv_std_logic_vector(6994,14),
		conv_std_logic_vector(6997,14),
		conv_std_logic_vector(7000,14),
		conv_std_logic_vector(7003,14),
		conv_std_logic_vector(7007,14),
		conv_std_logic_vector(7010,14),
		conv_std_logic_vector(7013,14),
		conv_std_logic_vector(7016,14),
		conv_std_logic_vector(7020,14),
		conv_std_logic_vector(7023,14),
		conv_std_logic_vector(7026,14),
		conv_std_logic_vector(7029,14),
		conv_std_logic_vector(7032,14),
		conv_std_logic_vector(7036,14),
		conv_std_logic_vector(7039,14),
		conv_std_logic_vector(7042,14),
		conv_std_logic_vector(7045,14),
		conv_std_logic_vector(7049,14),
		conv_std_logic_vector(7052,14),
		conv_std_logic_vector(7055,14),
		conv_std_logic_vector(7058,14),
		conv_std_logic_vector(7061,14),
		conv_std_logic_vector(7064,14),
		conv_std_logic_vector(7068,14),
		conv_std_logic_vector(7071,14),
		conv_std_logic_vector(7074,14),
		conv_std_logic_vector(7077,14),
		conv_std_logic_vector(7080,14),
		conv_std_logic_vector(7083,14),
		conv_std_logic_vector(7087,14),
		conv_std_logic_vector(7090,14),
		conv_std_logic_vector(7093,14),
		conv_std_logic_vector(7096,14),
		conv_std_logic_vector(7099,14),
		conv_std_logic_vector(7102,14),
		conv_std_logic_vector(7105,14),
		conv_std_logic_vector(7109,14),
		conv_std_logic_vector(7112,14),
		conv_std_logic_vector(7115,14),
		conv_std_logic_vector(7118,14),
		conv_std_logic_vector(7121,14),
		conv_std_logic_vector(7124,14),
		conv_std_logic_vector(7127,14),
		conv_std_logic_vector(7130,14),
		conv_std_logic_vector(7133,14),
		conv_std_logic_vector(7137,14),
		conv_std_logic_vector(7140,14),
		conv_std_logic_vector(7143,14),
		conv_std_logic_vector(7146,14),
		conv_std_logic_vector(7149,14),
		conv_std_logic_vector(7152,14),
		conv_std_logic_vector(7155,14),
		conv_std_logic_vector(7158,14),
		conv_std_logic_vector(7161,14),
		conv_std_logic_vector(7164,14),
		conv_std_logic_vector(7167,14),
		conv_std_logic_vector(7170,14),
		conv_std_logic_vector(7173,14),
		conv_std_logic_vector(7176,14),
		conv_std_logic_vector(7179,14),
		conv_std_logic_vector(7182,14),
		conv_std_logic_vector(7185,14),
		conv_std_logic_vector(7188,14),
		conv_std_logic_vector(7191,14),
		conv_std_logic_vector(7194,14),
		conv_std_logic_vector(7197,14),
		conv_std_logic_vector(7200,14),
		conv_std_logic_vector(7203,14),
		conv_std_logic_vector(7206,14),
		conv_std_logic_vector(7209,14),
		conv_std_logic_vector(7212,14),
		conv_std_logic_vector(7215,14),
		conv_std_logic_vector(7218,14),
		conv_std_logic_vector(7221,14),
		conv_std_logic_vector(7224,14),
		conv_std_logic_vector(7227,14),
		conv_std_logic_vector(7230,14),
		conv_std_logic_vector(7233,14),
		conv_std_logic_vector(7236,14),
		conv_std_logic_vector(7239,14),
		conv_std_logic_vector(7242,14),
		conv_std_logic_vector(7245,14),
		conv_std_logic_vector(7248,14),
		conv_std_logic_vector(7251,14),
		conv_std_logic_vector(7254,14),
		conv_std_logic_vector(7257,14),
		conv_std_logic_vector(7259,14),
		conv_std_logic_vector(7262,14),
		conv_std_logic_vector(7265,14),
		conv_std_logic_vector(7268,14),
		conv_std_logic_vector(7271,14),
		conv_std_logic_vector(7274,14),
		conv_std_logic_vector(7277,14),
		conv_std_logic_vector(7280,14),
		conv_std_logic_vector(7283,14),
		conv_std_logic_vector(7285,14),
		conv_std_logic_vector(7288,14),
		conv_std_logic_vector(7291,14),
		conv_std_logic_vector(7294,14),
		conv_std_logic_vector(7297,14),
		conv_std_logic_vector(7300,14),
		conv_std_logic_vector(7303,14),
		conv_std_logic_vector(7305,14),
		conv_std_logic_vector(7308,14),
		conv_std_logic_vector(7311,14),
		conv_std_logic_vector(7314,14),
		conv_std_logic_vector(7317,14),
		conv_std_logic_vector(7320,14),
		conv_std_logic_vector(7322,14),
		conv_std_logic_vector(7325,14),
		conv_std_logic_vector(7328,14),
		conv_std_logic_vector(7331,14),
		conv_std_logic_vector(7334,14),
		conv_std_logic_vector(7336,14),
		conv_std_logic_vector(7339,14),
		conv_std_logic_vector(7342,14),
		conv_std_logic_vector(7345,14),
		conv_std_logic_vector(7348,14),
		conv_std_logic_vector(7350,14),
		conv_std_logic_vector(7353,14),
		conv_std_logic_vector(7356,14),
		conv_std_logic_vector(7359,14),
		conv_std_logic_vector(7361,14),
		conv_std_logic_vector(7364,14),
		conv_std_logic_vector(7367,14),
		conv_std_logic_vector(7370,14),
		conv_std_logic_vector(7372,14),
		conv_std_logic_vector(7375,14),
		conv_std_logic_vector(7378,14),
		conv_std_logic_vector(7381,14),
		conv_std_logic_vector(7383,14),
		conv_std_logic_vector(7386,14),
		conv_std_logic_vector(7389,14),
		conv_std_logic_vector(7391,14),
		conv_std_logic_vector(7394,14),
		conv_std_logic_vector(7397,14),
		conv_std_logic_vector(7400,14),
		conv_std_logic_vector(7402,14),
		conv_std_logic_vector(7405,14),
		conv_std_logic_vector(7408,14),
		conv_std_logic_vector(7410,14),
		conv_std_logic_vector(7413,14),
		conv_std_logic_vector(7416,14),
		conv_std_logic_vector(7418,14),
		conv_std_logic_vector(7421,14),
		conv_std_logic_vector(7424,14),
		conv_std_logic_vector(7426,14),
		conv_std_logic_vector(7429,14),
		conv_std_logic_vector(7432,14),
		conv_std_logic_vector(7434,14),
		conv_std_logic_vector(7437,14),
		conv_std_logic_vector(7440,14),
		conv_std_logic_vector(7442,14),
		conv_std_logic_vector(7445,14),
		conv_std_logic_vector(7447,14),
		conv_std_logic_vector(7450,14),
		conv_std_logic_vector(7453,14),
		conv_std_logic_vector(7455,14),
		conv_std_logic_vector(7458,14),
		conv_std_logic_vector(7460,14),
		conv_std_logic_vector(7463,14),
		conv_std_logic_vector(7466,14),
		conv_std_logic_vector(7468,14),
		conv_std_logic_vector(7471,14),
		conv_std_logic_vector(7473,14),
		conv_std_logic_vector(7476,14),
		conv_std_logic_vector(7478,14),
		conv_std_logic_vector(7481,14),
		conv_std_logic_vector(7484,14),
		conv_std_logic_vector(7486,14),
		conv_std_logic_vector(7489,14),
		conv_std_logic_vector(7491,14),
		conv_std_logic_vector(7494,14),
		conv_std_logic_vector(7496,14),
		conv_std_logic_vector(7499,14),
		conv_std_logic_vector(7501,14),
		conv_std_logic_vector(7504,14),
		conv_std_logic_vector(7506,14),
		conv_std_logic_vector(7509,14),
		conv_std_logic_vector(7511,14),
		conv_std_logic_vector(7514,14),
		conv_std_logic_vector(7516,14),
		conv_std_logic_vector(7519,14),
		conv_std_logic_vector(7521,14),
		conv_std_logic_vector(7524,14),
		conv_std_logic_vector(7526,14),
		conv_std_logic_vector(7529,14),
		conv_std_logic_vector(7531,14),
		conv_std_logic_vector(7534,14),
		conv_std_logic_vector(7536,14),
		conv_std_logic_vector(7539,14),
		conv_std_logic_vector(7541,14),
		conv_std_logic_vector(7544,14),
		conv_std_logic_vector(7546,14),
		conv_std_logic_vector(7549,14),
		conv_std_logic_vector(7551,14),
		conv_std_logic_vector(7553,14),
		conv_std_logic_vector(7556,14),
		conv_std_logic_vector(7558,14),
		conv_std_logic_vector(7561,14),
		conv_std_logic_vector(7563,14),
		conv_std_logic_vector(7566,14),
		conv_std_logic_vector(7568,14),
		conv_std_logic_vector(7570,14),
		conv_std_logic_vector(7573,14),
		conv_std_logic_vector(7575,14),
		conv_std_logic_vector(7578,14),
		conv_std_logic_vector(7580,14),
		conv_std_logic_vector(7582,14),
		conv_std_logic_vector(7585,14),
		conv_std_logic_vector(7587,14),
		conv_std_logic_vector(7589,14),
		conv_std_logic_vector(7592,14),
		conv_std_logic_vector(7594,14),
		conv_std_logic_vector(7596,14),
		conv_std_logic_vector(7599,14),
		conv_std_logic_vector(7601,14),
		conv_std_logic_vector(7603,14),
		conv_std_logic_vector(7606,14),
		conv_std_logic_vector(7608,14),
		conv_std_logic_vector(7610,14),
		conv_std_logic_vector(7613,14),
		conv_std_logic_vector(7615,14),
		conv_std_logic_vector(7617,14),
		conv_std_logic_vector(7620,14),
		conv_std_logic_vector(7622,14),
		conv_std_logic_vector(7624,14),
		conv_std_logic_vector(7627,14),
		conv_std_logic_vector(7629,14),
		conv_std_logic_vector(7631,14),
		conv_std_logic_vector(7633,14),
		conv_std_logic_vector(7636,14),
		conv_std_logic_vector(7638,14),
		conv_std_logic_vector(7640,14),
		conv_std_logic_vector(7643,14),
		conv_std_logic_vector(7645,14),
		conv_std_logic_vector(7647,14),
		conv_std_logic_vector(7649,14),
		conv_std_logic_vector(7652,14),
		conv_std_logic_vector(7654,14),
		conv_std_logic_vector(7656,14),
		conv_std_logic_vector(7658,14),
		conv_std_logic_vector(7661,14),
		conv_std_logic_vector(7663,14),
		conv_std_logic_vector(7665,14),
		conv_std_logic_vector(7667,14),
		conv_std_logic_vector(7669,14),
		conv_std_logic_vector(7672,14),
		conv_std_logic_vector(7674,14),
		conv_std_logic_vector(7676,14),
		conv_std_logic_vector(7678,14),
		conv_std_logic_vector(7680,14),
		conv_std_logic_vector(7683,14),
		conv_std_logic_vector(7685,14),
		conv_std_logic_vector(7687,14),
		conv_std_logic_vector(7689,14),
		conv_std_logic_vector(7691,14),
		conv_std_logic_vector(7693,14),
		conv_std_logic_vector(7696,14),
		conv_std_logic_vector(7698,14),
		conv_std_logic_vector(7700,14),
		conv_std_logic_vector(7702,14),
		conv_std_logic_vector(7704,14),
		conv_std_logic_vector(7706,14),
		conv_std_logic_vector(7708,14),
		conv_std_logic_vector(7711,14),
		conv_std_logic_vector(7713,14),
		conv_std_logic_vector(7715,14),
		conv_std_logic_vector(7717,14),
		conv_std_logic_vector(7719,14),
		conv_std_logic_vector(7721,14),
		conv_std_logic_vector(7723,14),
		conv_std_logic_vector(7725,14),
		conv_std_logic_vector(7727,14),
		conv_std_logic_vector(7729,14),
		conv_std_logic_vector(7731,14),
		conv_std_logic_vector(7734,14),
		conv_std_logic_vector(7736,14),
		conv_std_logic_vector(7738,14),
		conv_std_logic_vector(7740,14),
		conv_std_logic_vector(7742,14),
		conv_std_logic_vector(7744,14),
		conv_std_logic_vector(7746,14),
		conv_std_logic_vector(7748,14),
		conv_std_logic_vector(7750,14),
		conv_std_logic_vector(7752,14),
		conv_std_logic_vector(7754,14),
		conv_std_logic_vector(7756,14),
		conv_std_logic_vector(7758,14),
		conv_std_logic_vector(7760,14),
		conv_std_logic_vector(7762,14),
		conv_std_logic_vector(7764,14),
		conv_std_logic_vector(7766,14),
		conv_std_logic_vector(7768,14),
		conv_std_logic_vector(7770,14),
		conv_std_logic_vector(7772,14),
		conv_std_logic_vector(7774,14),
		conv_std_logic_vector(7776,14),
		conv_std_logic_vector(7778,14),
		conv_std_logic_vector(7780,14),
		conv_std_logic_vector(7782,14),
		conv_std_logic_vector(7784,14),
		conv_std_logic_vector(7786,14),
		conv_std_logic_vector(7788,14),
		conv_std_logic_vector(7790,14),
		conv_std_logic_vector(7792,14),
		conv_std_logic_vector(7794,14),
		conv_std_logic_vector(7796,14),
		conv_std_logic_vector(7798,14),
		conv_std_logic_vector(7799,14),
		conv_std_logic_vector(7801,14),
		conv_std_logic_vector(7803,14),
		conv_std_logic_vector(7805,14),
		conv_std_logic_vector(7807,14),
		conv_std_logic_vector(7809,14),
		conv_std_logic_vector(7811,14),
		conv_std_logic_vector(7813,14),
		conv_std_logic_vector(7815,14),
		conv_std_logic_vector(7817,14),
		conv_std_logic_vector(7818,14),
		conv_std_logic_vector(7820,14),
		conv_std_logic_vector(7822,14),
		conv_std_logic_vector(7824,14),
		conv_std_logic_vector(7826,14),
		conv_std_logic_vector(7828,14),
		conv_std_logic_vector(7830,14),
		conv_std_logic_vector(7831,14),
		conv_std_logic_vector(7833,14),
		conv_std_logic_vector(7835,14),
		conv_std_logic_vector(7837,14),
		conv_std_logic_vector(7839,14),
		conv_std_logic_vector(7841,14),
		conv_std_logic_vector(7842,14),
		conv_std_logic_vector(7844,14),
		conv_std_logic_vector(7846,14),
		conv_std_logic_vector(7848,14),
		conv_std_logic_vector(7850,14),
		conv_std_logic_vector(7851,14),
		conv_std_logic_vector(7853,14),
		conv_std_logic_vector(7855,14),
		conv_std_logic_vector(7857,14),
		conv_std_logic_vector(7859,14),
		conv_std_logic_vector(7860,14),
		conv_std_logic_vector(7862,14),
		conv_std_logic_vector(7864,14),
		conv_std_logic_vector(7866,14),
		conv_std_logic_vector(7867,14),
		conv_std_logic_vector(7869,14),
		conv_std_logic_vector(7871,14),
		conv_std_logic_vector(7873,14),
		conv_std_logic_vector(7874,14),
		conv_std_logic_vector(7876,14),
		conv_std_logic_vector(7878,14),
		conv_std_logic_vector(7879,14),
		conv_std_logic_vector(7881,14),
		conv_std_logic_vector(7883,14),
		conv_std_logic_vector(7885,14),
		conv_std_logic_vector(7886,14),
		conv_std_logic_vector(7888,14),
		conv_std_logic_vector(7890,14),
		conv_std_logic_vector(7891,14),
		conv_std_logic_vector(7893,14),
		conv_std_logic_vector(7895,14),
		conv_std_logic_vector(7896,14),
		conv_std_logic_vector(7898,14),
		conv_std_logic_vector(7900,14),
		conv_std_logic_vector(7901,14),
		conv_std_logic_vector(7903,14),
		conv_std_logic_vector(7905,14),
		conv_std_logic_vector(7906,14),
		conv_std_logic_vector(7908,14),
		conv_std_logic_vector(7910,14),
		conv_std_logic_vector(7911,14),
		conv_std_logic_vector(7913,14),
		conv_std_logic_vector(7915,14),
		conv_std_logic_vector(7916,14),
		conv_std_logic_vector(7918,14),
		conv_std_logic_vector(7919,14),
		conv_std_logic_vector(7921,14),
		conv_std_logic_vector(7923,14),
		conv_std_logic_vector(7924,14),
		conv_std_logic_vector(7926,14),
		conv_std_logic_vector(7927,14),
		conv_std_logic_vector(7929,14),
		conv_std_logic_vector(7930,14),
		conv_std_logic_vector(7932,14),
		conv_std_logic_vector(7934,14),
		conv_std_logic_vector(7935,14),
		conv_std_logic_vector(7937,14),
		conv_std_logic_vector(7938,14),
		conv_std_logic_vector(7940,14),
		conv_std_logic_vector(7941,14),
		conv_std_logic_vector(7943,14),
		conv_std_logic_vector(7944,14),
		conv_std_logic_vector(7946,14),
		conv_std_logic_vector(7948,14),
		conv_std_logic_vector(7949,14),
		conv_std_logic_vector(7951,14),
		conv_std_logic_vector(7952,14),
		conv_std_logic_vector(7954,14),
		conv_std_logic_vector(7955,14),
		conv_std_logic_vector(7957,14),
		conv_std_logic_vector(7958,14),
		conv_std_logic_vector(7960,14),
		conv_std_logic_vector(7961,14),
		conv_std_logic_vector(7963,14),
		conv_std_logic_vector(7964,14),
		conv_std_logic_vector(7965,14),
		conv_std_logic_vector(7967,14),
		conv_std_logic_vector(7968,14),
		conv_std_logic_vector(7970,14),
		conv_std_logic_vector(7971,14),
		conv_std_logic_vector(7973,14),
		conv_std_logic_vector(7974,14),
		conv_std_logic_vector(7976,14),
		conv_std_logic_vector(7977,14),
		conv_std_logic_vector(7978,14),
		conv_std_logic_vector(7980,14),
		conv_std_logic_vector(7981,14),
		conv_std_logic_vector(7983,14),
		conv_std_logic_vector(7984,14),
		conv_std_logic_vector(7986,14),
		conv_std_logic_vector(7987,14),
		conv_std_logic_vector(7988,14),
		conv_std_logic_vector(7990,14),
		conv_std_logic_vector(7991,14),
		conv_std_logic_vector(7992,14),
		conv_std_logic_vector(7994,14),
		conv_std_logic_vector(7995,14),
		conv_std_logic_vector(7997,14),
		conv_std_logic_vector(7998,14),
		conv_std_logic_vector(7999,14),
		conv_std_logic_vector(8001,14),
		conv_std_logic_vector(8002,14),
		conv_std_logic_vector(8003,14),
		conv_std_logic_vector(8005,14),
		conv_std_logic_vector(8006,14),
		conv_std_logic_vector(8007,14),
		conv_std_logic_vector(8009,14),
		conv_std_logic_vector(8010,14),
		conv_std_logic_vector(8011,14),
		conv_std_logic_vector(8013,14),
		conv_std_logic_vector(8014,14),
		conv_std_logic_vector(8015,14),
		conv_std_logic_vector(8016,14),
		conv_std_logic_vector(8018,14),
		conv_std_logic_vector(8019,14),
		conv_std_logic_vector(8020,14),
		conv_std_logic_vector(8022,14),
		conv_std_logic_vector(8023,14),
		conv_std_logic_vector(8024,14),
		conv_std_logic_vector(8025,14),
		conv_std_logic_vector(8027,14),
		conv_std_logic_vector(8028,14),
		conv_std_logic_vector(8029,14),
		conv_std_logic_vector(8030,14),
		conv_std_logic_vector(8032,14),
		conv_std_logic_vector(8033,14),
		conv_std_logic_vector(8034,14),
		conv_std_logic_vector(8035,14),
		conv_std_logic_vector(8037,14),
		conv_std_logic_vector(8038,14),
		conv_std_logic_vector(8039,14),
		conv_std_logic_vector(8040,14),
		conv_std_logic_vector(8041,14),
		conv_std_logic_vector(8043,14),
		conv_std_logic_vector(8044,14),
		conv_std_logic_vector(8045,14),
		conv_std_logic_vector(8046,14),
		conv_std_logic_vector(8047,14),
		conv_std_logic_vector(8048,14),
		conv_std_logic_vector(8050,14),
		conv_std_logic_vector(8051,14),
		conv_std_logic_vector(8052,14),
		conv_std_logic_vector(8053,14),
		conv_std_logic_vector(8054,14),
		conv_std_logic_vector(8055,14),
		conv_std_logic_vector(8057,14),
		conv_std_logic_vector(8058,14),
		conv_std_logic_vector(8059,14),
		conv_std_logic_vector(8060,14),
		conv_std_logic_vector(8061,14),
		conv_std_logic_vector(8062,14),
		conv_std_logic_vector(8063,14),
		conv_std_logic_vector(8064,14),
		conv_std_logic_vector(8065,14),
		conv_std_logic_vector(8067,14),
		conv_std_logic_vector(8068,14),
		conv_std_logic_vector(8069,14),
		conv_std_logic_vector(8070,14),
		conv_std_logic_vector(8071,14),
		conv_std_logic_vector(8072,14),
		conv_std_logic_vector(8073,14),
		conv_std_logic_vector(8074,14),
		conv_std_logic_vector(8075,14),
		conv_std_logic_vector(8076,14),
		conv_std_logic_vector(8077,14),
		conv_std_logic_vector(8078,14),
		conv_std_logic_vector(8079,14),
		conv_std_logic_vector(8080,14),
		conv_std_logic_vector(8081,14),
		conv_std_logic_vector(8082,14),
		conv_std_logic_vector(8083,14),
		conv_std_logic_vector(8084,14),
		conv_std_logic_vector(8085,14),
		conv_std_logic_vector(8086,14),
		conv_std_logic_vector(8087,14),
		conv_std_logic_vector(8088,14),
		conv_std_logic_vector(8089,14),
		conv_std_logic_vector(8090,14),
		conv_std_logic_vector(8091,14),
		conv_std_logic_vector(8092,14),
		conv_std_logic_vector(8093,14),
		conv_std_logic_vector(8094,14),
		conv_std_logic_vector(8095,14),
		conv_std_logic_vector(8096,14),
		conv_std_logic_vector(8097,14),
		conv_std_logic_vector(8098,14),
		conv_std_logic_vector(8099,14),
		conv_std_logic_vector(8100,14),
		conv_std_logic_vector(8101,14),
		conv_std_logic_vector(8102,14),
		conv_std_logic_vector(8103,14),
		conv_std_logic_vector(8104,14),
		conv_std_logic_vector(8105,14),
		conv_std_logic_vector(8106,14),
		conv_std_logic_vector(8106,14),
		conv_std_logic_vector(8107,14),
		conv_std_logic_vector(8108,14),
		conv_std_logic_vector(8109,14),
		conv_std_logic_vector(8110,14),
		conv_std_logic_vector(8111,14),
		conv_std_logic_vector(8112,14),
		conv_std_logic_vector(8113,14),
		conv_std_logic_vector(8114,14),
		conv_std_logic_vector(8114,14),
		conv_std_logic_vector(8115,14),
		conv_std_logic_vector(8116,14),
		conv_std_logic_vector(8117,14),
		conv_std_logic_vector(8118,14),
		conv_std_logic_vector(8119,14),
		conv_std_logic_vector(8119,14),
		conv_std_logic_vector(8120,14),
		conv_std_logic_vector(8121,14),
		conv_std_logic_vector(8122,14),
		conv_std_logic_vector(8123,14),
		conv_std_logic_vector(8124,14),
		conv_std_logic_vector(8124,14),
		conv_std_logic_vector(8125,14),
		conv_std_logic_vector(8126,14),
		conv_std_logic_vector(8127,14),
		conv_std_logic_vector(8128,14),
		conv_std_logic_vector(8128,14),
		conv_std_logic_vector(8129,14),
		conv_std_logic_vector(8130,14),
		conv_std_logic_vector(8131,14),
		conv_std_logic_vector(8131,14),
		conv_std_logic_vector(8132,14),
		conv_std_logic_vector(8133,14),
		conv_std_logic_vector(8134,14),
		conv_std_logic_vector(8134,14),
		conv_std_logic_vector(8135,14),
		conv_std_logic_vector(8136,14),
		conv_std_logic_vector(8137,14),
		conv_std_logic_vector(8137,14),
		conv_std_logic_vector(8138,14),
		conv_std_logic_vector(8139,14),
		conv_std_logic_vector(8139,14),
		conv_std_logic_vector(8140,14),
		conv_std_logic_vector(8141,14),
		conv_std_logic_vector(8142,14),
		conv_std_logic_vector(8142,14),
		conv_std_logic_vector(8143,14),
		conv_std_logic_vector(8144,14),
		conv_std_logic_vector(8144,14),
		conv_std_logic_vector(8145,14),
		conv_std_logic_vector(8146,14),
		conv_std_logic_vector(8146,14),
		conv_std_logic_vector(8147,14),
		conv_std_logic_vector(8148,14),
		conv_std_logic_vector(8148,14),
		conv_std_logic_vector(8149,14),
		conv_std_logic_vector(8150,14),
		conv_std_logic_vector(8150,14),
		conv_std_logic_vector(8151,14),
		conv_std_logic_vector(8151,14),
		conv_std_logic_vector(8152,14),
		conv_std_logic_vector(8153,14),
		conv_std_logic_vector(8153,14),
		conv_std_logic_vector(8154,14),
		conv_std_logic_vector(8154,14),
		conv_std_logic_vector(8155,14),
		conv_std_logic_vector(8156,14),
		conv_std_logic_vector(8156,14),
		conv_std_logic_vector(8157,14),
		conv_std_logic_vector(8157,14),
		conv_std_logic_vector(8158,14),
		conv_std_logic_vector(8159,14),
		conv_std_logic_vector(8159,14),
		conv_std_logic_vector(8160,14),
		conv_std_logic_vector(8160,14),
		conv_std_logic_vector(8161,14),
		conv_std_logic_vector(8161,14),
		conv_std_logic_vector(8162,14),
		conv_std_logic_vector(8162,14),
		conv_std_logic_vector(8163,14),
		conv_std_logic_vector(8163,14),
		conv_std_logic_vector(8164,14),
		conv_std_logic_vector(8164,14),
		conv_std_logic_vector(8165,14),
		conv_std_logic_vector(8165,14),
		conv_std_logic_vector(8166,14),
		conv_std_logic_vector(8166,14),
		conv_std_logic_vector(8167,14),
		conv_std_logic_vector(8167,14),
		conv_std_logic_vector(8168,14),
		conv_std_logic_vector(8168,14),
		conv_std_logic_vector(8169,14),
		conv_std_logic_vector(8169,14),
		conv_std_logic_vector(8170,14),
		conv_std_logic_vector(8170,14),
		conv_std_logic_vector(8171,14),
		conv_std_logic_vector(8171,14),
		conv_std_logic_vector(8172,14),
		conv_std_logic_vector(8172,14),
		conv_std_logic_vector(8172,14),
		conv_std_logic_vector(8173,14),
		conv_std_logic_vector(8173,14),
		conv_std_logic_vector(8174,14),
		conv_std_logic_vector(8174,14),
		conv_std_logic_vector(8175,14),
		conv_std_logic_vector(8175,14),
		conv_std_logic_vector(8175,14),
		conv_std_logic_vector(8176,14),
		conv_std_logic_vector(8176,14),
		conv_std_logic_vector(8176,14),
		conv_std_logic_vector(8177,14),
		conv_std_logic_vector(8177,14),
		conv_std_logic_vector(8178,14),
		conv_std_logic_vector(8178,14),
		conv_std_logic_vector(8178,14),
		conv_std_logic_vector(8179,14),
		conv_std_logic_vector(8179,14),
		conv_std_logic_vector(8179,14),
		conv_std_logic_vector(8180,14),
		conv_std_logic_vector(8180,14),
		conv_std_logic_vector(8180,14),
		conv_std_logic_vector(8181,14),
		conv_std_logic_vector(8181,14),
		conv_std_logic_vector(8181,14),
		conv_std_logic_vector(8182,14),
		conv_std_logic_vector(8182,14),
		conv_std_logic_vector(8182,14),
		conv_std_logic_vector(8183,14),
		conv_std_logic_vector(8183,14),
		conv_std_logic_vector(8183,14),
		conv_std_logic_vector(8183,14),
		conv_std_logic_vector(8184,14),
		conv_std_logic_vector(8184,14),
		conv_std_logic_vector(8184,14),
		conv_std_logic_vector(8184,14),
		conv_std_logic_vector(8185,14),
		conv_std_logic_vector(8185,14),
		conv_std_logic_vector(8185,14),
		conv_std_logic_vector(8185,14),
		conv_std_logic_vector(8186,14),
		conv_std_logic_vector(8186,14),
		conv_std_logic_vector(8186,14),
		conv_std_logic_vector(8186,14),
		conv_std_logic_vector(8187,14),
		conv_std_logic_vector(8187,14),
		conv_std_logic_vector(8187,14),
		conv_std_logic_vector(8187,14),
		conv_std_logic_vector(8187,14),
		conv_std_logic_vector(8188,14),
		conv_std_logic_vector(8188,14),
		conv_std_logic_vector(8188,14),
		conv_std_logic_vector(8188,14),
		conv_std_logic_vector(8188,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8192,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8191,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8190,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8189,14),
		conv_std_logic_vector(8188,14),
		conv_std_logic_vector(8188,14),
		conv_std_logic_vector(8188,14),
		conv_std_logic_vector(8188,14),
		conv_std_logic_vector(8188,14),
		conv_std_logic_vector(8187,14),
		conv_std_logic_vector(8187,14),
		conv_std_logic_vector(8187,14),
		conv_std_logic_vector(8187,14),
		conv_std_logic_vector(8187,14),
		conv_std_logic_vector(8186,14),
		conv_std_logic_vector(8186,14),
		conv_std_logic_vector(8186,14),
		conv_std_logic_vector(8186,14),
		conv_std_logic_vector(8185,14),
		conv_std_logic_vector(8185,14),
		conv_std_logic_vector(8185,14),
		conv_std_logic_vector(8185,14),
		conv_std_logic_vector(8184,14),
		conv_std_logic_vector(8184,14),
		conv_std_logic_vector(8184,14),
		conv_std_logic_vector(8184,14),
		conv_std_logic_vector(8183,14),
		conv_std_logic_vector(8183,14),
		conv_std_logic_vector(8183,14),
		conv_std_logic_vector(8183,14),
		conv_std_logic_vector(8182,14),
		conv_std_logic_vector(8182,14),
		conv_std_logic_vector(8182,14),
		conv_std_logic_vector(8181,14),
		conv_std_logic_vector(8181,14),
		conv_std_logic_vector(8181,14),
		conv_std_logic_vector(8180,14),
		conv_std_logic_vector(8180,14),
		conv_std_logic_vector(8180,14),
		conv_std_logic_vector(8179,14),
		conv_std_logic_vector(8179,14),
		conv_std_logic_vector(8179,14),
		conv_std_logic_vector(8178,14),
		conv_std_logic_vector(8178,14),
		conv_std_logic_vector(8178,14),
		conv_std_logic_vector(8177,14),
		conv_std_logic_vector(8177,14),
		conv_std_logic_vector(8176,14),
		conv_std_logic_vector(8176,14),
		conv_std_logic_vector(8176,14),
		conv_std_logic_vector(8175,14),
		conv_std_logic_vector(8175,14),
		conv_std_logic_vector(8175,14),
		conv_std_logic_vector(8174,14),
		conv_std_logic_vector(8174,14),
		conv_std_logic_vector(8173,14),
		conv_std_logic_vector(8173,14),
		conv_std_logic_vector(8172,14),
		conv_std_logic_vector(8172,14),
		conv_std_logic_vector(8172,14),
		conv_std_logic_vector(8171,14),
		conv_std_logic_vector(8171,14),
		conv_std_logic_vector(8170,14),
		conv_std_logic_vector(8170,14),
		conv_std_logic_vector(8169,14),
		conv_std_logic_vector(8169,14),
		conv_std_logic_vector(8168,14),
		conv_std_logic_vector(8168,14),
		conv_std_logic_vector(8167,14),
		conv_std_logic_vector(8167,14),
		conv_std_logic_vector(8166,14),
		conv_std_logic_vector(8166,14),
		conv_std_logic_vector(8165,14),
		conv_std_logic_vector(8165,14),
		conv_std_logic_vector(8164,14),
		conv_std_logic_vector(8164,14),
		conv_std_logic_vector(8163,14),
		conv_std_logic_vector(8163,14),
		conv_std_logic_vector(8162,14),
		conv_std_logic_vector(8162,14),
		conv_std_logic_vector(8161,14),
		conv_std_logic_vector(8161,14),
		conv_std_logic_vector(8160,14),
		conv_std_logic_vector(8160,14),
		conv_std_logic_vector(8159,14),
		conv_std_logic_vector(8159,14),
		conv_std_logic_vector(8158,14),
		conv_std_logic_vector(8157,14),
		conv_std_logic_vector(8157,14),
		conv_std_logic_vector(8156,14),
		conv_std_logic_vector(8156,14),
		conv_std_logic_vector(8155,14),
		conv_std_logic_vector(8154,14),
		conv_std_logic_vector(8154,14),
		conv_std_logic_vector(8153,14),
		conv_std_logic_vector(8153,14),
		conv_std_logic_vector(8152,14),
		conv_std_logic_vector(8151,14),
		conv_std_logic_vector(8151,14),
		conv_std_logic_vector(8150,14),
		conv_std_logic_vector(8150,14),
		conv_std_logic_vector(8149,14),
		conv_std_logic_vector(8148,14),
		conv_std_logic_vector(8148,14),
		conv_std_logic_vector(8147,14),
		conv_std_logic_vector(8146,14),
		conv_std_logic_vector(8146,14),
		conv_std_logic_vector(8145,14),
		conv_std_logic_vector(8144,14),
		conv_std_logic_vector(8144,14),
		conv_std_logic_vector(8143,14),
		conv_std_logic_vector(8142,14),
		conv_std_logic_vector(8142,14),
		conv_std_logic_vector(8141,14),
		conv_std_logic_vector(8140,14),
		conv_std_logic_vector(8139,14),
		conv_std_logic_vector(8139,14),
		conv_std_logic_vector(8138,14),
		conv_std_logic_vector(8137,14),
		conv_std_logic_vector(8137,14),
		conv_std_logic_vector(8136,14),
		conv_std_logic_vector(8135,14),
		conv_std_logic_vector(8134,14),
		conv_std_logic_vector(8134,14),
		conv_std_logic_vector(8133,14),
		conv_std_logic_vector(8132,14),
		conv_std_logic_vector(8131,14),
		conv_std_logic_vector(8131,14),
		conv_std_logic_vector(8130,14),
		conv_std_logic_vector(8129,14),
		conv_std_logic_vector(8128,14),
		conv_std_logic_vector(8128,14),
		conv_std_logic_vector(8127,14),
		conv_std_logic_vector(8126,14),
		conv_std_logic_vector(8125,14),
		conv_std_logic_vector(8124,14),
		conv_std_logic_vector(8124,14),
		conv_std_logic_vector(8123,14),
		conv_std_logic_vector(8122,14),
		conv_std_logic_vector(8121,14),
		conv_std_logic_vector(8120,14),
		conv_std_logic_vector(8119,14),
		conv_std_logic_vector(8119,14),
		conv_std_logic_vector(8118,14),
		conv_std_logic_vector(8117,14),
		conv_std_logic_vector(8116,14),
		conv_std_logic_vector(8115,14),
		conv_std_logic_vector(8114,14),
		conv_std_logic_vector(8114,14),
		conv_std_logic_vector(8113,14),
		conv_std_logic_vector(8112,14),
		conv_std_logic_vector(8111,14),
		conv_std_logic_vector(8110,14),
		conv_std_logic_vector(8109,14),
		conv_std_logic_vector(8108,14),
		conv_std_logic_vector(8107,14),
		conv_std_logic_vector(8106,14),
		conv_std_logic_vector(8106,14),
		conv_std_logic_vector(8105,14),
		conv_std_logic_vector(8104,14),
		conv_std_logic_vector(8103,14),
		conv_std_logic_vector(8102,14),
		conv_std_logic_vector(8101,14),
		conv_std_logic_vector(8100,14),
		conv_std_logic_vector(8099,14),
		conv_std_logic_vector(8098,14),
		conv_std_logic_vector(8097,14),
		conv_std_logic_vector(8096,14),
		conv_std_logic_vector(8095,14),
		conv_std_logic_vector(8094,14),
		conv_std_logic_vector(8093,14),
		conv_std_logic_vector(8092,14),
		conv_std_logic_vector(8091,14),
		conv_std_logic_vector(8090,14),
		conv_std_logic_vector(8089,14),
		conv_std_logic_vector(8088,14),
		conv_std_logic_vector(8087,14),
		conv_std_logic_vector(8086,14),
		conv_std_logic_vector(8085,14),
		conv_std_logic_vector(8084,14),
		conv_std_logic_vector(8083,14),
		conv_std_logic_vector(8082,14),
		conv_std_logic_vector(8081,14),
		conv_std_logic_vector(8080,14),
		conv_std_logic_vector(8079,14),
		conv_std_logic_vector(8078,14),
		conv_std_logic_vector(8077,14),
		conv_std_logic_vector(8076,14),
		conv_std_logic_vector(8075,14),
		conv_std_logic_vector(8074,14),
		conv_std_logic_vector(8073,14),
		conv_std_logic_vector(8072,14),
		conv_std_logic_vector(8071,14),
		conv_std_logic_vector(8070,14),
		conv_std_logic_vector(8069,14),
		conv_std_logic_vector(8068,14),
		conv_std_logic_vector(8067,14),
		conv_std_logic_vector(8065,14),
		conv_std_logic_vector(8064,14),
		conv_std_logic_vector(8063,14),
		conv_std_logic_vector(8062,14),
		conv_std_logic_vector(8061,14),
		conv_std_logic_vector(8060,14),
		conv_std_logic_vector(8059,14),
		conv_std_logic_vector(8058,14),
		conv_std_logic_vector(8057,14),
		conv_std_logic_vector(8055,14),
		conv_std_logic_vector(8054,14),
		conv_std_logic_vector(8053,14),
		conv_std_logic_vector(8052,14),
		conv_std_logic_vector(8051,14),
		conv_std_logic_vector(8050,14),
		conv_std_logic_vector(8048,14),
		conv_std_logic_vector(8047,14),
		conv_std_logic_vector(8046,14),
		conv_std_logic_vector(8045,14),
		conv_std_logic_vector(8044,14),
		conv_std_logic_vector(8043,14),
		conv_std_logic_vector(8041,14),
		conv_std_logic_vector(8040,14),
		conv_std_logic_vector(8039,14),
		conv_std_logic_vector(8038,14),
		conv_std_logic_vector(8037,14),
		conv_std_logic_vector(8035,14),
		conv_std_logic_vector(8034,14),
		conv_std_logic_vector(8033,14),
		conv_std_logic_vector(8032,14),
		conv_std_logic_vector(8030,14),
		conv_std_logic_vector(8029,14),
		conv_std_logic_vector(8028,14),
		conv_std_logic_vector(8027,14),
		conv_std_logic_vector(8025,14),
		conv_std_logic_vector(8024,14),
		conv_std_logic_vector(8023,14),
		conv_std_logic_vector(8022,14),
		conv_std_logic_vector(8020,14),
		conv_std_logic_vector(8019,14),
		conv_std_logic_vector(8018,14),
		conv_std_logic_vector(8016,14),
		conv_std_logic_vector(8015,14),
		conv_std_logic_vector(8014,14),
		conv_std_logic_vector(8013,14),
		conv_std_logic_vector(8011,14),
		conv_std_logic_vector(8010,14),
		conv_std_logic_vector(8009,14),
		conv_std_logic_vector(8007,14),
		conv_std_logic_vector(8006,14),
		conv_std_logic_vector(8005,14),
		conv_std_logic_vector(8003,14),
		conv_std_logic_vector(8002,14),
		conv_std_logic_vector(8001,14),
		conv_std_logic_vector(7999,14),
		conv_std_logic_vector(7998,14),
		conv_std_logic_vector(7997,14),
		conv_std_logic_vector(7995,14),
		conv_std_logic_vector(7994,14),
		conv_std_logic_vector(7992,14),
		conv_std_logic_vector(7991,14),
		conv_std_logic_vector(7990,14),
		conv_std_logic_vector(7988,14),
		conv_std_logic_vector(7987,14),
		conv_std_logic_vector(7986,14),
		conv_std_logic_vector(7984,14),
		conv_std_logic_vector(7983,14),
		conv_std_logic_vector(7981,14),
		conv_std_logic_vector(7980,14),
		conv_std_logic_vector(7978,14),
		conv_std_logic_vector(7977,14),
		conv_std_logic_vector(7976,14),
		conv_std_logic_vector(7974,14),
		conv_std_logic_vector(7973,14),
		conv_std_logic_vector(7971,14),
		conv_std_logic_vector(7970,14),
		conv_std_logic_vector(7968,14),
		conv_std_logic_vector(7967,14),
		conv_std_logic_vector(7965,14),
		conv_std_logic_vector(7964,14),
		conv_std_logic_vector(7963,14),
		conv_std_logic_vector(7961,14),
		conv_std_logic_vector(7960,14),
		conv_std_logic_vector(7958,14),
		conv_std_logic_vector(7957,14),
		conv_std_logic_vector(7955,14),
		conv_std_logic_vector(7954,14),
		conv_std_logic_vector(7952,14),
		conv_std_logic_vector(7951,14),
		conv_std_logic_vector(7949,14),
		conv_std_logic_vector(7948,14),
		conv_std_logic_vector(7946,14),
		conv_std_logic_vector(7944,14),
		conv_std_logic_vector(7943,14),
		conv_std_logic_vector(7941,14),
		conv_std_logic_vector(7940,14),
		conv_std_logic_vector(7938,14),
		conv_std_logic_vector(7937,14),
		conv_std_logic_vector(7935,14),
		conv_std_logic_vector(7934,14),
		conv_std_logic_vector(7932,14),
		conv_std_logic_vector(7930,14),
		conv_std_logic_vector(7929,14),
		conv_std_logic_vector(7927,14),
		conv_std_logic_vector(7926,14),
		conv_std_logic_vector(7924,14),
		conv_std_logic_vector(7923,14),
		conv_std_logic_vector(7921,14),
		conv_std_logic_vector(7919,14),
		conv_std_logic_vector(7918,14),
		conv_std_logic_vector(7916,14),
		conv_std_logic_vector(7915,14),
		conv_std_logic_vector(7913,14),
		conv_std_logic_vector(7911,14),
		conv_std_logic_vector(7910,14),
		conv_std_logic_vector(7908,14),
		conv_std_logic_vector(7906,14),
		conv_std_logic_vector(7905,14),
		conv_std_logic_vector(7903,14),
		conv_std_logic_vector(7901,14),
		conv_std_logic_vector(7900,14),
		conv_std_logic_vector(7898,14),
		conv_std_logic_vector(7896,14),
		conv_std_logic_vector(7895,14),
		conv_std_logic_vector(7893,14),
		conv_std_logic_vector(7891,14),
		conv_std_logic_vector(7890,14),
		conv_std_logic_vector(7888,14),
		conv_std_logic_vector(7886,14),
		conv_std_logic_vector(7885,14),
		conv_std_logic_vector(7883,14),
		conv_std_logic_vector(7881,14),
		conv_std_logic_vector(7879,14),
		conv_std_logic_vector(7878,14),
		conv_std_logic_vector(7876,14),
		conv_std_logic_vector(7874,14),
		conv_std_logic_vector(7873,14),
		conv_std_logic_vector(7871,14),
		conv_std_logic_vector(7869,14),
		conv_std_logic_vector(7867,14),
		conv_std_logic_vector(7866,14),
		conv_std_logic_vector(7864,14),
		conv_std_logic_vector(7862,14),
		conv_std_logic_vector(7860,14),
		conv_std_logic_vector(7859,14),
		conv_std_logic_vector(7857,14),
		conv_std_logic_vector(7855,14),
		conv_std_logic_vector(7853,14),
		conv_std_logic_vector(7851,14),
		conv_std_logic_vector(7850,14),
		conv_std_logic_vector(7848,14),
		conv_std_logic_vector(7846,14),
		conv_std_logic_vector(7844,14),
		conv_std_logic_vector(7842,14),
		conv_std_logic_vector(7841,14),
		conv_std_logic_vector(7839,14),
		conv_std_logic_vector(7837,14),
		conv_std_logic_vector(7835,14),
		conv_std_logic_vector(7833,14),
		conv_std_logic_vector(7831,14),
		conv_std_logic_vector(7830,14),
		conv_std_logic_vector(7828,14),
		conv_std_logic_vector(7826,14),
		conv_std_logic_vector(7824,14),
		conv_std_logic_vector(7822,14),
		conv_std_logic_vector(7820,14),
		conv_std_logic_vector(7818,14),
		conv_std_logic_vector(7817,14),
		conv_std_logic_vector(7815,14),
		conv_std_logic_vector(7813,14),
		conv_std_logic_vector(7811,14),
		conv_std_logic_vector(7809,14),
		conv_std_logic_vector(7807,14),
		conv_std_logic_vector(7805,14),
		conv_std_logic_vector(7803,14),
		conv_std_logic_vector(7801,14),
		conv_std_logic_vector(7799,14),
		conv_std_logic_vector(7798,14),
		conv_std_logic_vector(7796,14),
		conv_std_logic_vector(7794,14),
		conv_std_logic_vector(7792,14),
		conv_std_logic_vector(7790,14),
		conv_std_logic_vector(7788,14),
		conv_std_logic_vector(7786,14),
		conv_std_logic_vector(7784,14),
		conv_std_logic_vector(7782,14),
		conv_std_logic_vector(7780,14),
		conv_std_logic_vector(7778,14),
		conv_std_logic_vector(7776,14),
		conv_std_logic_vector(7774,14),
		conv_std_logic_vector(7772,14),
		conv_std_logic_vector(7770,14),
		conv_std_logic_vector(7768,14),
		conv_std_logic_vector(7766,14),
		conv_std_logic_vector(7764,14),
		conv_std_logic_vector(7762,14),
		conv_std_logic_vector(7760,14),
		conv_std_logic_vector(7758,14),
		conv_std_logic_vector(7756,14),
		conv_std_logic_vector(7754,14),
		conv_std_logic_vector(7752,14),
		conv_std_logic_vector(7750,14),
		conv_std_logic_vector(7748,14),
		conv_std_logic_vector(7746,14),
		conv_std_logic_vector(7744,14),
		conv_std_logic_vector(7742,14),
		conv_std_logic_vector(7740,14),
		conv_std_logic_vector(7738,14),
		conv_std_logic_vector(7736,14),
		conv_std_logic_vector(7734,14),
		conv_std_logic_vector(7731,14),
		conv_std_logic_vector(7729,14),
		conv_std_logic_vector(7727,14),
		conv_std_logic_vector(7725,14),
		conv_std_logic_vector(7723,14),
		conv_std_logic_vector(7721,14),
		conv_std_logic_vector(7719,14),
		conv_std_logic_vector(7717,14),
		conv_std_logic_vector(7715,14),
		conv_std_logic_vector(7713,14),
		conv_std_logic_vector(7711,14),
		conv_std_logic_vector(7708,14),
		conv_std_logic_vector(7706,14),
		conv_std_logic_vector(7704,14),
		conv_std_logic_vector(7702,14),
		conv_std_logic_vector(7700,14),
		conv_std_logic_vector(7698,14),
		conv_std_logic_vector(7696,14),
		conv_std_logic_vector(7693,14),
		conv_std_logic_vector(7691,14),
		conv_std_logic_vector(7689,14),
		conv_std_logic_vector(7687,14),
		conv_std_logic_vector(7685,14),
		conv_std_logic_vector(7683,14),
		conv_std_logic_vector(7680,14),
		conv_std_logic_vector(7678,14),
		conv_std_logic_vector(7676,14),
		conv_std_logic_vector(7674,14),
		conv_std_logic_vector(7672,14),
		conv_std_logic_vector(7669,14),
		conv_std_logic_vector(7667,14),
		conv_std_logic_vector(7665,14),
		conv_std_logic_vector(7663,14),
		conv_std_logic_vector(7661,14),
		conv_std_logic_vector(7658,14),
		conv_std_logic_vector(7656,14),
		conv_std_logic_vector(7654,14),
		conv_std_logic_vector(7652,14),
		conv_std_logic_vector(7649,14),
		conv_std_logic_vector(7647,14),
		conv_std_logic_vector(7645,14),
		conv_std_logic_vector(7643,14),
		conv_std_logic_vector(7640,14),
		conv_std_logic_vector(7638,14),
		conv_std_logic_vector(7636,14),
		conv_std_logic_vector(7633,14),
		conv_std_logic_vector(7631,14),
		conv_std_logic_vector(7629,14),
		conv_std_logic_vector(7627,14),
		conv_std_logic_vector(7624,14),
		conv_std_logic_vector(7622,14),
		conv_std_logic_vector(7620,14),
		conv_std_logic_vector(7617,14),
		conv_std_logic_vector(7615,14),
		conv_std_logic_vector(7613,14),
		conv_std_logic_vector(7610,14),
		conv_std_logic_vector(7608,14),
		conv_std_logic_vector(7606,14),
		conv_std_logic_vector(7603,14),
		conv_std_logic_vector(7601,14),
		conv_std_logic_vector(7599,14),
		conv_std_logic_vector(7596,14),
		conv_std_logic_vector(7594,14),
		conv_std_logic_vector(7592,14),
		conv_std_logic_vector(7589,14),
		conv_std_logic_vector(7587,14),
		conv_std_logic_vector(7585,14),
		conv_std_logic_vector(7582,14),
		conv_std_logic_vector(7580,14),
		conv_std_logic_vector(7578,14),
		conv_std_logic_vector(7575,14),
		conv_std_logic_vector(7573,14),
		conv_std_logic_vector(7570,14),
		conv_std_logic_vector(7568,14),
		conv_std_logic_vector(7566,14),
		conv_std_logic_vector(7563,14),
		conv_std_logic_vector(7561,14),
		conv_std_logic_vector(7558,14),
		conv_std_logic_vector(7556,14),
		conv_std_logic_vector(7553,14),
		conv_std_logic_vector(7551,14),
		conv_std_logic_vector(7549,14),
		conv_std_logic_vector(7546,14),
		conv_std_logic_vector(7544,14),
		conv_std_logic_vector(7541,14),
		conv_std_logic_vector(7539,14),
		conv_std_logic_vector(7536,14),
		conv_std_logic_vector(7534,14),
		conv_std_logic_vector(7531,14),
		conv_std_logic_vector(7529,14),
		conv_std_logic_vector(7526,14),
		conv_std_logic_vector(7524,14),
		conv_std_logic_vector(7521,14),
		conv_std_logic_vector(7519,14),
		conv_std_logic_vector(7516,14),
		conv_std_logic_vector(7514,14),
		conv_std_logic_vector(7511,14),
		conv_std_logic_vector(7509,14),
		conv_std_logic_vector(7506,14),
		conv_std_logic_vector(7504,14),
		conv_std_logic_vector(7501,14),
		conv_std_logic_vector(7499,14),
		conv_std_logic_vector(7496,14),
		conv_std_logic_vector(7494,14),
		conv_std_logic_vector(7491,14),
		conv_std_logic_vector(7489,14),
		conv_std_logic_vector(7486,14),
		conv_std_logic_vector(7484,14),
		conv_std_logic_vector(7481,14),
		conv_std_logic_vector(7478,14),
		conv_std_logic_vector(7476,14),
		conv_std_logic_vector(7473,14),
		conv_std_logic_vector(7471,14),
		conv_std_logic_vector(7468,14),
		conv_std_logic_vector(7466,14),
		conv_std_logic_vector(7463,14),
		conv_std_logic_vector(7460,14),
		conv_std_logic_vector(7458,14),
		conv_std_logic_vector(7455,14),
		conv_std_logic_vector(7453,14),
		conv_std_logic_vector(7450,14),
		conv_std_logic_vector(7447,14),
		conv_std_logic_vector(7445,14),
		conv_std_logic_vector(7442,14),
		conv_std_logic_vector(7440,14),
		conv_std_logic_vector(7437,14),
		conv_std_logic_vector(7434,14),
		conv_std_logic_vector(7432,14),
		conv_std_logic_vector(7429,14),
		conv_std_logic_vector(7426,14),
		conv_std_logic_vector(7424,14),
		conv_std_logic_vector(7421,14),
		conv_std_logic_vector(7418,14),
		conv_std_logic_vector(7416,14),
		conv_std_logic_vector(7413,14),
		conv_std_logic_vector(7410,14),
		conv_std_logic_vector(7408,14),
		conv_std_logic_vector(7405,14),
		conv_std_logic_vector(7402,14),
		conv_std_logic_vector(7400,14),
		conv_std_logic_vector(7397,14),
		conv_std_logic_vector(7394,14),
		conv_std_logic_vector(7391,14),
		conv_std_logic_vector(7389,14),
		conv_std_logic_vector(7386,14),
		conv_std_logic_vector(7383,14),
		conv_std_logic_vector(7381,14),
		conv_std_logic_vector(7378,14),
		conv_std_logic_vector(7375,14),
		conv_std_logic_vector(7372,14),
		conv_std_logic_vector(7370,14),
		conv_std_logic_vector(7367,14),
		conv_std_logic_vector(7364,14),
		conv_std_logic_vector(7361,14),
		conv_std_logic_vector(7359,14),
		conv_std_logic_vector(7356,14),
		conv_std_logic_vector(7353,14),
		conv_std_logic_vector(7350,14),
		conv_std_logic_vector(7348,14),
		conv_std_logic_vector(7345,14),
		conv_std_logic_vector(7342,14),
		conv_std_logic_vector(7339,14),
		conv_std_logic_vector(7336,14),
		conv_std_logic_vector(7334,14),
		conv_std_logic_vector(7331,14),
		conv_std_logic_vector(7328,14),
		conv_std_logic_vector(7325,14),
		conv_std_logic_vector(7322,14),
		conv_std_logic_vector(7320,14),
		conv_std_logic_vector(7317,14),
		conv_std_logic_vector(7314,14),
		conv_std_logic_vector(7311,14),
		conv_std_logic_vector(7308,14),
		conv_std_logic_vector(7305,14),
		conv_std_logic_vector(7303,14),
		conv_std_logic_vector(7300,14),
		conv_std_logic_vector(7297,14),
		conv_std_logic_vector(7294,14),
		conv_std_logic_vector(7291,14),
		conv_std_logic_vector(7288,14),
		conv_std_logic_vector(7285,14),
		conv_std_logic_vector(7283,14),
		conv_std_logic_vector(7280,14),
		conv_std_logic_vector(7277,14),
		conv_std_logic_vector(7274,14),
		conv_std_logic_vector(7271,14),
		conv_std_logic_vector(7268,14),
		conv_std_logic_vector(7265,14),
		conv_std_logic_vector(7262,14),
		conv_std_logic_vector(7259,14),
		conv_std_logic_vector(7257,14),
		conv_std_logic_vector(7254,14),
		conv_std_logic_vector(7251,14),
		conv_std_logic_vector(7248,14),
		conv_std_logic_vector(7245,14),
		conv_std_logic_vector(7242,14),
		conv_std_logic_vector(7239,14),
		conv_std_logic_vector(7236,14),
		conv_std_logic_vector(7233,14),
		conv_std_logic_vector(7230,14),
		conv_std_logic_vector(7227,14),
		conv_std_logic_vector(7224,14),
		conv_std_logic_vector(7221,14),
		conv_std_logic_vector(7218,14),
		conv_std_logic_vector(7215,14),
		conv_std_logic_vector(7212,14),
		conv_std_logic_vector(7209,14),
		conv_std_logic_vector(7206,14),
		conv_std_logic_vector(7203,14),
		conv_std_logic_vector(7200,14),
		conv_std_logic_vector(7197,14),
		conv_std_logic_vector(7194,14),
		conv_std_logic_vector(7191,14),
		conv_std_logic_vector(7188,14),
		conv_std_logic_vector(7185,14),
		conv_std_logic_vector(7182,14),
		conv_std_logic_vector(7179,14),
		conv_std_logic_vector(7176,14),
		conv_std_logic_vector(7173,14),
		conv_std_logic_vector(7170,14),
		conv_std_logic_vector(7167,14),
		conv_std_logic_vector(7164,14),
		conv_std_logic_vector(7161,14),
		conv_std_logic_vector(7158,14),
		conv_std_logic_vector(7155,14),
		conv_std_logic_vector(7152,14),
		conv_std_logic_vector(7149,14),
		conv_std_logic_vector(7146,14),
		conv_std_logic_vector(7143,14),
		conv_std_logic_vector(7140,14),
		conv_std_logic_vector(7137,14),
		conv_std_logic_vector(7133,14),
		conv_std_logic_vector(7130,14),
		conv_std_logic_vector(7127,14),
		conv_std_logic_vector(7124,14),
		conv_std_logic_vector(7121,14),
		conv_std_logic_vector(7118,14),
		conv_std_logic_vector(7115,14),
		conv_std_logic_vector(7112,14),
		conv_std_logic_vector(7109,14),
		conv_std_logic_vector(7105,14),
		conv_std_logic_vector(7102,14),
		conv_std_logic_vector(7099,14),
		conv_std_logic_vector(7096,14),
		conv_std_logic_vector(7093,14),
		conv_std_logic_vector(7090,14),
		conv_std_logic_vector(7087,14),
		conv_std_logic_vector(7083,14),
		conv_std_logic_vector(7080,14),
		conv_std_logic_vector(7077,14),
		conv_std_logic_vector(7074,14),
		conv_std_logic_vector(7071,14),
		conv_std_logic_vector(7068,14),
		conv_std_logic_vector(7064,14),
		conv_std_logic_vector(7061,14),
		conv_std_logic_vector(7058,14),
		conv_std_logic_vector(7055,14),
		conv_std_logic_vector(7052,14),
		conv_std_logic_vector(7049,14),
		conv_std_logic_vector(7045,14),
		conv_std_logic_vector(7042,14),
		conv_std_logic_vector(7039,14),
		conv_std_logic_vector(7036,14),
		conv_std_logic_vector(7032,14),
		conv_std_logic_vector(7029,14),
		conv_std_logic_vector(7026,14),
		conv_std_logic_vector(7023,14),
		conv_std_logic_vector(7020,14),
		conv_std_logic_vector(7016,14),
		conv_std_logic_vector(7013,14),
		conv_std_logic_vector(7010,14),
		conv_std_logic_vector(7007,14),
		conv_std_logic_vector(7003,14),
		conv_std_logic_vector(7000,14),
		conv_std_logic_vector(6997,14),
		conv_std_logic_vector(6994,14),
		conv_std_logic_vector(6990,14),
		conv_std_logic_vector(6987,14),
		conv_std_logic_vector(6984,14),
		conv_std_logic_vector(6980,14),
		conv_std_logic_vector(6977,14),
		conv_std_logic_vector(6974,14),
		conv_std_logic_vector(6971,14),
		conv_std_logic_vector(6967,14),
		conv_std_logic_vector(6964,14),
		conv_std_logic_vector(6961,14),
		conv_std_logic_vector(6957,14),
		conv_std_logic_vector(6954,14),
		conv_std_logic_vector(6951,14),
		conv_std_logic_vector(6947,14),
		conv_std_logic_vector(6944,14),
		conv_std_logic_vector(6941,14),
		conv_std_logic_vector(6937,14),
		conv_std_logic_vector(6934,14),
		conv_std_logic_vector(6931,14),
		conv_std_logic_vector(6927,14),
		conv_std_logic_vector(6924,14),
		conv_std_logic_vector(6921,14),
		conv_std_logic_vector(6917,14),
		conv_std_logic_vector(6914,14),
		conv_std_logic_vector(6910,14),
		conv_std_logic_vector(6907,14),
		conv_std_logic_vector(6904,14),
		conv_std_logic_vector(6900,14),
		conv_std_logic_vector(6897,14),
		conv_std_logic_vector(6894,14),
		conv_std_logic_vector(6890,14),
		conv_std_logic_vector(6887,14),
		conv_std_logic_vector(6883,14),
		conv_std_logic_vector(6880,14),
		conv_std_logic_vector(6876,14),
		conv_std_logic_vector(6873,14),
		conv_std_logic_vector(6870,14),
		conv_std_logic_vector(6866,14),
		conv_std_logic_vector(6863,14),
		conv_std_logic_vector(6859,14),
		conv_std_logic_vector(6856,14),
		conv_std_logic_vector(6852,14),
		conv_std_logic_vector(6849,14),
		conv_std_logic_vector(6846,14),
		conv_std_logic_vector(6842,14),
		conv_std_logic_vector(6839,14),
		conv_std_logic_vector(6835,14),
		conv_std_logic_vector(6832,14),
		conv_std_logic_vector(6828,14),
		conv_std_logic_vector(6825,14),
		conv_std_logic_vector(6821,14),
		conv_std_logic_vector(6818,14),
		conv_std_logic_vector(6814,14),
		conv_std_logic_vector(6811,14),
		conv_std_logic_vector(6807,14),
		conv_std_logic_vector(6804,14),
		conv_std_logic_vector(6800,14),
		conv_std_logic_vector(6797,14),
		conv_std_logic_vector(6793,14),
		conv_std_logic_vector(6790,14),
		conv_std_logic_vector(6786,14),
		conv_std_logic_vector(6783,14),
		conv_std_logic_vector(6779,14),
		conv_std_logic_vector(6776,14),
		conv_std_logic_vector(6772,14),
		conv_std_logic_vector(6769,14),
		conv_std_logic_vector(6765,14),
		conv_std_logic_vector(6762,14),
		conv_std_logic_vector(6758,14),
		conv_std_logic_vector(6755,14),
		conv_std_logic_vector(6751,14),
		conv_std_logic_vector(6747,14),
		conv_std_logic_vector(6744,14),
		conv_std_logic_vector(6740,14),
		conv_std_logic_vector(6737,14),
		conv_std_logic_vector(6733,14),
		conv_std_logic_vector(6730,14),
		conv_std_logic_vector(6726,14),
		conv_std_logic_vector(6722,14),
		conv_std_logic_vector(6719,14),
		conv_std_logic_vector(6715,14),
		conv_std_logic_vector(6712,14),
		conv_std_logic_vector(6708,14),
		conv_std_logic_vector(6704,14),
		conv_std_logic_vector(6701,14),
		conv_std_logic_vector(6697,14),
		conv_std_logic_vector(6694,14),
		conv_std_logic_vector(6690,14),
		conv_std_logic_vector(6686,14),
		conv_std_logic_vector(6683,14),
		conv_std_logic_vector(6679,14),
		conv_std_logic_vector(6675,14),
		conv_std_logic_vector(6672,14),
		conv_std_logic_vector(6668,14),
		conv_std_logic_vector(6664,14),
		conv_std_logic_vector(6661,14),
		conv_std_logic_vector(6657,14),
		conv_std_logic_vector(6653,14),
		conv_std_logic_vector(6650,14),
		conv_std_logic_vector(6646,14),
		conv_std_logic_vector(6642,14),
		conv_std_logic_vector(6639,14),
		conv_std_logic_vector(6635,14),
		conv_std_logic_vector(6631,14),
		conv_std_logic_vector(6628,14),
		conv_std_logic_vector(6624,14),
		conv_std_logic_vector(6620,14),
		conv_std_logic_vector(6617,14),
		conv_std_logic_vector(6613,14),
		conv_std_logic_vector(6609,14),
		conv_std_logic_vector(6605,14),
		conv_std_logic_vector(6602,14),
		conv_std_logic_vector(6598,14),
		conv_std_logic_vector(6594,14),
		conv_std_logic_vector(6591,14),
		conv_std_logic_vector(6587,14),
		conv_std_logic_vector(6583,14),
		conv_std_logic_vector(6579,14),
		conv_std_logic_vector(6576,14),
		conv_std_logic_vector(6572,14),
		conv_std_logic_vector(6568,14),
		conv_std_logic_vector(6564,14),
		conv_std_logic_vector(6561,14),
		conv_std_logic_vector(6557,14),
		conv_std_logic_vector(6553,14),
		conv_std_logic_vector(6549,14),
		conv_std_logic_vector(6546,14),
		conv_std_logic_vector(6542,14),
		conv_std_logic_vector(6538,14),
		conv_std_logic_vector(6534,14),
		conv_std_logic_vector(6530,14),
		conv_std_logic_vector(6527,14),
		conv_std_logic_vector(6523,14),
		conv_std_logic_vector(6519,14),
		conv_std_logic_vector(6515,14),
		conv_std_logic_vector(6511,14),
		conv_std_logic_vector(6508,14),
		conv_std_logic_vector(6504,14),
		conv_std_logic_vector(6500,14),
		conv_std_logic_vector(6496,14),
		conv_std_logic_vector(6492,14),
		conv_std_logic_vector(6488,14),
		conv_std_logic_vector(6485,14),
		conv_std_logic_vector(6481,14),
		conv_std_logic_vector(6477,14),
		conv_std_logic_vector(6473,14),
		conv_std_logic_vector(6469,14),
		conv_std_logic_vector(6465,14),
		conv_std_logic_vector(6461,14),
		conv_std_logic_vector(6458,14),
		conv_std_logic_vector(6454,14),
		conv_std_logic_vector(6450,14),
		conv_std_logic_vector(6446,14),
		conv_std_logic_vector(6442,14),
		conv_std_logic_vector(6438,14),
		conv_std_logic_vector(6434,14),
		conv_std_logic_vector(6430,14),
		conv_std_logic_vector(6427,14),
		conv_std_logic_vector(6423,14),
		conv_std_logic_vector(6419,14),
		conv_std_logic_vector(6415,14),
		conv_std_logic_vector(6411,14),
		conv_std_logic_vector(6407,14),
		conv_std_logic_vector(6403,14),
		conv_std_logic_vector(6399,14),
		conv_std_logic_vector(6395,14),
		conv_std_logic_vector(6391,14),
		conv_std_logic_vector(6387,14),
		conv_std_logic_vector(6384,14),
		conv_std_logic_vector(6380,14),
		conv_std_logic_vector(6376,14),
		conv_std_logic_vector(6372,14),
		conv_std_logic_vector(6368,14),
		conv_std_logic_vector(6364,14),
		conv_std_logic_vector(6360,14),
		conv_std_logic_vector(6356,14),
		conv_std_logic_vector(6352,14),
		conv_std_logic_vector(6348,14),
		conv_std_logic_vector(6344,14),
		conv_std_logic_vector(6340,14),
		conv_std_logic_vector(6336,14),
		conv_std_logic_vector(6332,14),
		conv_std_logic_vector(6328,14),
		conv_std_logic_vector(6324,14),
		conv_std_logic_vector(6320,14),
		conv_std_logic_vector(6316,14),
		conv_std_logic_vector(6312,14),
		conv_std_logic_vector(6308,14),
		conv_std_logic_vector(6304,14),
		conv_std_logic_vector(6300,14),
		conv_std_logic_vector(6296,14),
		conv_std_logic_vector(6292,14),
		conv_std_logic_vector(6288,14),
		conv_std_logic_vector(6284,14),
		conv_std_logic_vector(6280,14),
		conv_std_logic_vector(6276,14),
		conv_std_logic_vector(6272,14),
		conv_std_logic_vector(6268,14),
		conv_std_logic_vector(6264,14),
		conv_std_logic_vector(6260,14),
		conv_std_logic_vector(6256,14),
		conv_std_logic_vector(6252,14),
		conv_std_logic_vector(6247,14),
		conv_std_logic_vector(6243,14),
		conv_std_logic_vector(6239,14),
		conv_std_logic_vector(6235,14),
		conv_std_logic_vector(6231,14),
		conv_std_logic_vector(6227,14),
		conv_std_logic_vector(6223,14),
		conv_std_logic_vector(6219,14),
		conv_std_logic_vector(6215,14),
		conv_std_logic_vector(6211,14),
		conv_std_logic_vector(6207,14),
		conv_std_logic_vector(6203,14),
		conv_std_logic_vector(6198,14),
		conv_std_logic_vector(6194,14),
		conv_std_logic_vector(6190,14),
		conv_std_logic_vector(6186,14),
		conv_std_logic_vector(6182,14),
		conv_std_logic_vector(6178,14),
		conv_std_logic_vector(6174,14),
		conv_std_logic_vector(6170,14),
		conv_std_logic_vector(6165,14),
		conv_std_logic_vector(6161,14),
		conv_std_logic_vector(6157,14),
		conv_std_logic_vector(6153,14),
		conv_std_logic_vector(6149,14),
		conv_std_logic_vector(6145,14),
		conv_std_logic_vector(6141,14),
		conv_std_logic_vector(6136,14),
		conv_std_logic_vector(6132,14),
		conv_std_logic_vector(6128,14),
		conv_std_logic_vector(6124,14),
		conv_std_logic_vector(6120,14),
		conv_std_logic_vector(6116,14),
		conv_std_logic_vector(6111,14),
		conv_std_logic_vector(6107,14),
		conv_std_logic_vector(6103,14),
		conv_std_logic_vector(6099,14),
		conv_std_logic_vector(6095,14),
		conv_std_logic_vector(6090,14),
		conv_std_logic_vector(6086,14),
		conv_std_logic_vector(6082,14),
		conv_std_logic_vector(6078,14),
		conv_std_logic_vector(6074,14),
		conv_std_logic_vector(6069,14),
		conv_std_logic_vector(6065,14),
		conv_std_logic_vector(6061,14),
		conv_std_logic_vector(6057,14),
		conv_std_logic_vector(6052,14),
		conv_std_logic_vector(6048,14),
		conv_std_logic_vector(6044,14),
		conv_std_logic_vector(6040,14),
		conv_std_logic_vector(6036,14),
		conv_std_logic_vector(6031,14),
		conv_std_logic_vector(6027,14),
		conv_std_logic_vector(6023,14),
		conv_std_logic_vector(6018,14),
		conv_std_logic_vector(6014,14),
		conv_std_logic_vector(6010,14),
		conv_std_logic_vector(6006,14),
		conv_std_logic_vector(6001,14),
		conv_std_logic_vector(5997,14),
		conv_std_logic_vector(5993,14),
		conv_std_logic_vector(5989,14),
		conv_std_logic_vector(5984,14),
		conv_std_logic_vector(5980,14),
		conv_std_logic_vector(5976,14),
		conv_std_logic_vector(5971,14),
		conv_std_logic_vector(5967,14),
		conv_std_logic_vector(5963,14),
		conv_std_logic_vector(5958,14),
		conv_std_logic_vector(5954,14),
		conv_std_logic_vector(5950,14),
		conv_std_logic_vector(5946,14),
		conv_std_logic_vector(5941,14),
		conv_std_logic_vector(5937,14),
		conv_std_logic_vector(5933,14),
		conv_std_logic_vector(5928,14),
		conv_std_logic_vector(5924,14),
		conv_std_logic_vector(5920,14),
		conv_std_logic_vector(5915,14),
		conv_std_logic_vector(5911,14),
		conv_std_logic_vector(5906,14),
		conv_std_logic_vector(5902,14),
		conv_std_logic_vector(5898,14),
		conv_std_logic_vector(5893,14),
		conv_std_logic_vector(5889,14),
		conv_std_logic_vector(5885,14),
		conv_std_logic_vector(5880,14),
		conv_std_logic_vector(5876,14),
		conv_std_logic_vector(5872,14),
		conv_std_logic_vector(5867,14),
		conv_std_logic_vector(5863,14),
		conv_std_logic_vector(5858,14),
		conv_std_logic_vector(5854,14),
		conv_std_logic_vector(5850,14),
		conv_std_logic_vector(5845,14),
		conv_std_logic_vector(5841,14),
		conv_std_logic_vector(5836,14),
		conv_std_logic_vector(5832,14),
		conv_std_logic_vector(5828,14),
		conv_std_logic_vector(5823,14),
		conv_std_logic_vector(5819,14),
		conv_std_logic_vector(5814,14),
		conv_std_logic_vector(5810,14),
		conv_std_logic_vector(5805,14),
		conv_std_logic_vector(5801,14),
		conv_std_logic_vector(5797,14),
		conv_std_logic_vector(5792,14),
		conv_std_logic_vector(5788,14),
		conv_std_logic_vector(5783,14),
		conv_std_logic_vector(5779,14),
		conv_std_logic_vector(5774,14),
		conv_std_logic_vector(5770,14),
		conv_std_logic_vector(5765,14),
		conv_std_logic_vector(5761,14),
		conv_std_logic_vector(5756,14),
		conv_std_logic_vector(5752,14),
		conv_std_logic_vector(5748,14),
		conv_std_logic_vector(5743,14),
		conv_std_logic_vector(5739,14),
		conv_std_logic_vector(5734,14),
		conv_std_logic_vector(5730,14),
		conv_std_logic_vector(5725,14),
		conv_std_logic_vector(5721,14),
		conv_std_logic_vector(5716,14),
		conv_std_logic_vector(5712,14),
		conv_std_logic_vector(5707,14),
		conv_std_logic_vector(5703,14),
		conv_std_logic_vector(5698,14),
		conv_std_logic_vector(5694,14),
		conv_std_logic_vector(5689,14),
		conv_std_logic_vector(5685,14),
		conv_std_logic_vector(5680,14),
		conv_std_logic_vector(5675,14),
		conv_std_logic_vector(5671,14),
		conv_std_logic_vector(5666,14),
		conv_std_logic_vector(5662,14),
		conv_std_logic_vector(5657,14),
		conv_std_logic_vector(5653,14),
		conv_std_logic_vector(5648,14),
		conv_std_logic_vector(5644,14),
		conv_std_logic_vector(5639,14),
		conv_std_logic_vector(5635,14),
		conv_std_logic_vector(5630,14),
		conv_std_logic_vector(5625,14),
		conv_std_logic_vector(5621,14),
		conv_std_logic_vector(5616,14),
		conv_std_logic_vector(5612,14),
		conv_std_logic_vector(5607,14),
		conv_std_logic_vector(5603,14),
		conv_std_logic_vector(5598,14),
		conv_std_logic_vector(5593,14),
		conv_std_logic_vector(5589,14),
		conv_std_logic_vector(5584,14),
		conv_std_logic_vector(5580,14),
		conv_std_logic_vector(5575,14),
		conv_std_logic_vector(5570,14),
		conv_std_logic_vector(5566,14),
		conv_std_logic_vector(5561,14),
		conv_std_logic_vector(5557,14),
		conv_std_logic_vector(5552,14),
		conv_std_logic_vector(5547,14),
		conv_std_logic_vector(5543,14),
		conv_std_logic_vector(5538,14),
		conv_std_logic_vector(5533,14),
		conv_std_logic_vector(5529,14),
		conv_std_logic_vector(5524,14),
		conv_std_logic_vector(5520,14),
		conv_std_logic_vector(5515,14),
		conv_std_logic_vector(5510,14),
		conv_std_logic_vector(5506,14),
		conv_std_logic_vector(5501,14),
		conv_std_logic_vector(5496,14),
		conv_std_logic_vector(5492,14),
		conv_std_logic_vector(5487,14),
		conv_std_logic_vector(5482,14),
		conv_std_logic_vector(5478,14),
		conv_std_logic_vector(5473,14),
		conv_std_logic_vector(5468,14),
		conv_std_logic_vector(5464,14),
		conv_std_logic_vector(5459,14),
		conv_std_logic_vector(5454,14),
		conv_std_logic_vector(5450,14),
		conv_std_logic_vector(5445,14),
		conv_std_logic_vector(5440,14),
		conv_std_logic_vector(5435,14),
		conv_std_logic_vector(5431,14),
		conv_std_logic_vector(5426,14),
		conv_std_logic_vector(5421,14),
		conv_std_logic_vector(5417,14),
		conv_std_logic_vector(5412,14),
		conv_std_logic_vector(5407,14),
		conv_std_logic_vector(5402,14),
		conv_std_logic_vector(5398,14),
		conv_std_logic_vector(5393,14),
		conv_std_logic_vector(5388,14),
		conv_std_logic_vector(5384,14),
		conv_std_logic_vector(5379,14),
		conv_std_logic_vector(5374,14),
		conv_std_logic_vector(5369,14),
		conv_std_logic_vector(5365,14),
		conv_std_logic_vector(5360,14),
		conv_std_logic_vector(5355,14),
		conv_std_logic_vector(5350,14),
		conv_std_logic_vector(5346,14),
		conv_std_logic_vector(5341,14),
		conv_std_logic_vector(5336,14),
		conv_std_logic_vector(5331,14),
		conv_std_logic_vector(5326,14),
		conv_std_logic_vector(5322,14),
		conv_std_logic_vector(5317,14),
		conv_std_logic_vector(5312,14),
		conv_std_logic_vector(5307,14),
		conv_std_logic_vector(5303,14),
		conv_std_logic_vector(5298,14),
		conv_std_logic_vector(5293,14),
		conv_std_logic_vector(5288,14),
		conv_std_logic_vector(5283,14),
		conv_std_logic_vector(5279,14),
		conv_std_logic_vector(5274,14),
		conv_std_logic_vector(5269,14),
		conv_std_logic_vector(5264,14),
		conv_std_logic_vector(5259,14),
		conv_std_logic_vector(5255,14),
		conv_std_logic_vector(5250,14),
		conv_std_logic_vector(5245,14),
		conv_std_logic_vector(5240,14),
		conv_std_logic_vector(5235,14),
		conv_std_logic_vector(5230,14),
		conv_std_logic_vector(5226,14),
		conv_std_logic_vector(5221,14),
		conv_std_logic_vector(5216,14),
		conv_std_logic_vector(5211,14),
		conv_std_logic_vector(5206,14),
		conv_std_logic_vector(5201,14),
		conv_std_logic_vector(5196,14),
		conv_std_logic_vector(5192,14),
		conv_std_logic_vector(5187,14),
		conv_std_logic_vector(5182,14),
		conv_std_logic_vector(5177,14),
		conv_std_logic_vector(5172,14),
		conv_std_logic_vector(5167,14),
		conv_std_logic_vector(5162,14),
		conv_std_logic_vector(5157,14),
		conv_std_logic_vector(5153,14),
		conv_std_logic_vector(5148,14),
		conv_std_logic_vector(5143,14),
		conv_std_logic_vector(5138,14),
		conv_std_logic_vector(5133,14),
		conv_std_logic_vector(5128,14),
		conv_std_logic_vector(5123,14),
		conv_std_logic_vector(5118,14),
		conv_std_logic_vector(5113,14),
		conv_std_logic_vector(5109,14),
		conv_std_logic_vector(5104,14),
		conv_std_logic_vector(5099,14),
		conv_std_logic_vector(5094,14),
		conv_std_logic_vector(5089,14),
		conv_std_logic_vector(5084,14),
		conv_std_logic_vector(5079,14),
		conv_std_logic_vector(5074,14),
		conv_std_logic_vector(5069,14),
		conv_std_logic_vector(5064,14),
		conv_std_logic_vector(5059,14),
		conv_std_logic_vector(5054,14),
		conv_std_logic_vector(5049,14),
		conv_std_logic_vector(5044,14),
		conv_std_logic_vector(5039,14),
		conv_std_logic_vector(5035,14),
		conv_std_logic_vector(5030,14),
		conv_std_logic_vector(5025,14),
		conv_std_logic_vector(5020,14),
		conv_std_logic_vector(5015,14),
		conv_std_logic_vector(5010,14),
		conv_std_logic_vector(5005,14),
		conv_std_logic_vector(5000,14),
		conv_std_logic_vector(4995,14),
		conv_std_logic_vector(4990,14),
		conv_std_logic_vector(4985,14),
		conv_std_logic_vector(4980,14),
		conv_std_logic_vector(4975,14),
		conv_std_logic_vector(4970,14),
		conv_std_logic_vector(4965,14),
		conv_std_logic_vector(4960,14),
		conv_std_logic_vector(4955,14),
		conv_std_logic_vector(4950,14),
		conv_std_logic_vector(4945,14),
		conv_std_logic_vector(4940,14),
		conv_std_logic_vector(4935,14),
		conv_std_logic_vector(4930,14),
		conv_std_logic_vector(4925,14),
		conv_std_logic_vector(4920,14),
		conv_std_logic_vector(4915,14),
		conv_std_logic_vector(4910,14),
		conv_std_logic_vector(4905,14),
		conv_std_logic_vector(4900,14),
		conv_std_logic_vector(4895,14),
		conv_std_logic_vector(4890,14),
		conv_std_logic_vector(4885,14),
		conv_std_logic_vector(4879,14),
		conv_std_logic_vector(4874,14),
		conv_std_logic_vector(4869,14),
		conv_std_logic_vector(4864,14),
		conv_std_logic_vector(4859,14),
		conv_std_logic_vector(4854,14),
		conv_std_logic_vector(4849,14),
		conv_std_logic_vector(4844,14),
		conv_std_logic_vector(4839,14),
		conv_std_logic_vector(4834,14),
		conv_std_logic_vector(4829,14),
		conv_std_logic_vector(4824,14),
		conv_std_logic_vector(4819,14),
		conv_std_logic_vector(4814,14),
		conv_std_logic_vector(4809,14),
		conv_std_logic_vector(4803,14),
		conv_std_logic_vector(4798,14),
		conv_std_logic_vector(4793,14),
		conv_std_logic_vector(4788,14),
		conv_std_logic_vector(4783,14),
		conv_std_logic_vector(4778,14),
		conv_std_logic_vector(4773,14),
		conv_std_logic_vector(4768,14),
		conv_std_logic_vector(4763,14),
		conv_std_logic_vector(4758,14),
		conv_std_logic_vector(4752,14),
		conv_std_logic_vector(4747,14),
		conv_std_logic_vector(4742,14),
		conv_std_logic_vector(4737,14),
		conv_std_logic_vector(4732,14),
		conv_std_logic_vector(4727,14),
		conv_std_logic_vector(4722,14),
		conv_std_logic_vector(4717,14),
		conv_std_logic_vector(4711,14),
		conv_std_logic_vector(4706,14),
		conv_std_logic_vector(4701,14),
		conv_std_logic_vector(4696,14),
		conv_std_logic_vector(4691,14),
		conv_std_logic_vector(4686,14),
		conv_std_logic_vector(4680,14),
		conv_std_logic_vector(4675,14),
		conv_std_logic_vector(4670,14),
		conv_std_logic_vector(4665,14),
		conv_std_logic_vector(4660,14),
		conv_std_logic_vector(4655,14),
		conv_std_logic_vector(4650,14),
		conv_std_logic_vector(4644,14),
		conv_std_logic_vector(4639,14),
		conv_std_logic_vector(4634,14),
		conv_std_logic_vector(4629,14),
		conv_std_logic_vector(4624,14),
		conv_std_logic_vector(4618,14),
		conv_std_logic_vector(4613,14),
		conv_std_logic_vector(4608,14),
		conv_std_logic_vector(4603,14),
		conv_std_logic_vector(4598,14),
		conv_std_logic_vector(4592,14),
		conv_std_logic_vector(4587,14),
		conv_std_logic_vector(4582,14),
		conv_std_logic_vector(4577,14),
		conv_std_logic_vector(4572,14),
		conv_std_logic_vector(4566,14),
		conv_std_logic_vector(4561,14),
		conv_std_logic_vector(4556,14),
		conv_std_logic_vector(4551,14),
		conv_std_logic_vector(4546,14),
		conv_std_logic_vector(4540,14),
		conv_std_logic_vector(4535,14),
		conv_std_logic_vector(4530,14),
		conv_std_logic_vector(4525,14),
		conv_std_logic_vector(4519,14),
		conv_std_logic_vector(4514,14),
		conv_std_logic_vector(4509,14),
		conv_std_logic_vector(4504,14),
		conv_std_logic_vector(4498,14),
		conv_std_logic_vector(4493,14),
		conv_std_logic_vector(4488,14),
		conv_std_logic_vector(4483,14),
		conv_std_logic_vector(4477,14),
		conv_std_logic_vector(4472,14),
		conv_std_logic_vector(4467,14),
		conv_std_logic_vector(4462,14),
		conv_std_logic_vector(4456,14),
		conv_std_logic_vector(4451,14),
		conv_std_logic_vector(4446,14),
		conv_std_logic_vector(4440,14),
		conv_std_logic_vector(4435,14),
		conv_std_logic_vector(4430,14),
		conv_std_logic_vector(4425,14),
		conv_std_logic_vector(4419,14),
		conv_std_logic_vector(4414,14),
		conv_std_logic_vector(4409,14),
		conv_std_logic_vector(4403,14),
		conv_std_logic_vector(4398,14),
		conv_std_logic_vector(4393,14),
		conv_std_logic_vector(4388,14),
		conv_std_logic_vector(4382,14),
		conv_std_logic_vector(4377,14),
		conv_std_logic_vector(4372,14),
		conv_std_logic_vector(4366,14),
		conv_std_logic_vector(4361,14),
		conv_std_logic_vector(4356,14),
		conv_std_logic_vector(4350,14),
		conv_std_logic_vector(4345,14),
		conv_std_logic_vector(4340,14),
		conv_std_logic_vector(4334,14),
		conv_std_logic_vector(4329,14),
		conv_std_logic_vector(4324,14),
		conv_std_logic_vector(4318,14),
		conv_std_logic_vector(4313,14),
		conv_std_logic_vector(4308,14),
		conv_std_logic_vector(4302,14),
		conv_std_logic_vector(4297,14),
		conv_std_logic_vector(4292,14),
		conv_std_logic_vector(4286,14),
		conv_std_logic_vector(4281,14),
		conv_std_logic_vector(4276,14),
		conv_std_logic_vector(4270,14),
		conv_std_logic_vector(4265,14),
		conv_std_logic_vector(4259,14),
		conv_std_logic_vector(4254,14),
		conv_std_logic_vector(4249,14),
		conv_std_logic_vector(4243,14),
		conv_std_logic_vector(4238,14),
		conv_std_logic_vector(4233,14),
		conv_std_logic_vector(4227,14),
		conv_std_logic_vector(4222,14),
		conv_std_logic_vector(4216,14),
		conv_std_logic_vector(4211,14),
		conv_std_logic_vector(4206,14),
		conv_std_logic_vector(4200,14),
		conv_std_logic_vector(4195,14),
		conv_std_logic_vector(4189,14),
		conv_std_logic_vector(4184,14),
		conv_std_logic_vector(4179,14),
		conv_std_logic_vector(4173,14),
		conv_std_logic_vector(4168,14),
		conv_std_logic_vector(4162,14),
		conv_std_logic_vector(4157,14),
		conv_std_logic_vector(4152,14),
		conv_std_logic_vector(4146,14),
		conv_std_logic_vector(4141,14),
		conv_std_logic_vector(4135,14),
		conv_std_logic_vector(4130,14),
		conv_std_logic_vector(4124,14),
		conv_std_logic_vector(4119,14),
		conv_std_logic_vector(4114,14),
		conv_std_logic_vector(4108,14),
		conv_std_logic_vector(4103,14),
		conv_std_logic_vector(4097,14),
		conv_std_logic_vector(4092,14),
		conv_std_logic_vector(4086,14),
		conv_std_logic_vector(4081,14),
		conv_std_logic_vector(4076,14),
		conv_std_logic_vector(4070,14),
		conv_std_logic_vector(4065,14),
		conv_std_logic_vector(4059,14),
		conv_std_logic_vector(4054,14),
		conv_std_logic_vector(4048,14),
		conv_std_logic_vector(4043,14),
		conv_std_logic_vector(4037,14),
		conv_std_logic_vector(4032,14),
		conv_std_logic_vector(4026,14),
		conv_std_logic_vector(4021,14),
		conv_std_logic_vector(4015,14),
		conv_std_logic_vector(4010,14),
		conv_std_logic_vector(4004,14),
		conv_std_logic_vector(3999,14),
		conv_std_logic_vector(3994,14),
		conv_std_logic_vector(3988,14),
		conv_std_logic_vector(3983,14),
		conv_std_logic_vector(3977,14),
		conv_std_logic_vector(3972,14),
		conv_std_logic_vector(3966,14),
		conv_std_logic_vector(3961,14),
		conv_std_logic_vector(3955,14),
		conv_std_logic_vector(3950,14),
		conv_std_logic_vector(3944,14),
		conv_std_logic_vector(3939,14),
		conv_std_logic_vector(3933,14),
		conv_std_logic_vector(3928,14),
		conv_std_logic_vector(3922,14),
		conv_std_logic_vector(3916,14),
		conv_std_logic_vector(3911,14),
		conv_std_logic_vector(3905,14),
		conv_std_logic_vector(3900,14),
		conv_std_logic_vector(3894,14),
		conv_std_logic_vector(3889,14),
		conv_std_logic_vector(3883,14),
		conv_std_logic_vector(3878,14),
		conv_std_logic_vector(3872,14),
		conv_std_logic_vector(3867,14),
		conv_std_logic_vector(3861,14),
		conv_std_logic_vector(3856,14),
		conv_std_logic_vector(3850,14),
		conv_std_logic_vector(3845,14),
		conv_std_logic_vector(3839,14),
		conv_std_logic_vector(3833,14),
		conv_std_logic_vector(3828,14),
		conv_std_logic_vector(3822,14),
		conv_std_logic_vector(3817,14),
		conv_std_logic_vector(3811,14),
		conv_std_logic_vector(3806,14),
		conv_std_logic_vector(3800,14),
		conv_std_logic_vector(3795,14),
		conv_std_logic_vector(3789,14),
		conv_std_logic_vector(3783,14),
		conv_std_logic_vector(3778,14),
		conv_std_logic_vector(3772,14),
		conv_std_logic_vector(3767,14),
		conv_std_logic_vector(3761,14),
		conv_std_logic_vector(3755,14),
		conv_std_logic_vector(3750,14),
		conv_std_logic_vector(3744,14),
		conv_std_logic_vector(3739,14),
		conv_std_logic_vector(3733,14),
		conv_std_logic_vector(3728,14),
		conv_std_logic_vector(3722,14),
		conv_std_logic_vector(3716,14),
		conv_std_logic_vector(3711,14),
		conv_std_logic_vector(3705,14),
		conv_std_logic_vector(3700,14),
		conv_std_logic_vector(3694,14),
		conv_std_logic_vector(3688,14),
		conv_std_logic_vector(3683,14),
		conv_std_logic_vector(3677,14),
		conv_std_logic_vector(3671,14),
		conv_std_logic_vector(3666,14),
		conv_std_logic_vector(3660,14),
		conv_std_logic_vector(3655,14),
		conv_std_logic_vector(3649,14),
		conv_std_logic_vector(3643,14),
		conv_std_logic_vector(3638,14),
		conv_std_logic_vector(3632,14),
		conv_std_logic_vector(3626,14),
		conv_std_logic_vector(3621,14),
		conv_std_logic_vector(3615,14),
		conv_std_logic_vector(3610,14),
		conv_std_logic_vector(3604,14),
		conv_std_logic_vector(3598,14),
		conv_std_logic_vector(3593,14),
		conv_std_logic_vector(3587,14),
		conv_std_logic_vector(3581,14),
		conv_std_logic_vector(3576,14),
		conv_std_logic_vector(3570,14),
		conv_std_logic_vector(3564,14),
		conv_std_logic_vector(3559,14),
		conv_std_logic_vector(3553,14),
		conv_std_logic_vector(3547,14),
		conv_std_logic_vector(3542,14),
		conv_std_logic_vector(3536,14),
		conv_std_logic_vector(3530,14),
		conv_std_logic_vector(3525,14),
		conv_std_logic_vector(3519,14),
		conv_std_logic_vector(3513,14),
		conv_std_logic_vector(3508,14),
		conv_std_logic_vector(3502,14),
		conv_std_logic_vector(3496,14),
		conv_std_logic_vector(3491,14),
		conv_std_logic_vector(3485,14),
		conv_std_logic_vector(3479,14),
		conv_std_logic_vector(3474,14),
		conv_std_logic_vector(3468,14),
		conv_std_logic_vector(3462,14),
		conv_std_logic_vector(3457,14),
		conv_std_logic_vector(3451,14),
		conv_std_logic_vector(3445,14),
		conv_std_logic_vector(3439,14),
		conv_std_logic_vector(3434,14),
		conv_std_logic_vector(3428,14),
		conv_std_logic_vector(3422,14),
		conv_std_logic_vector(3417,14),
		conv_std_logic_vector(3411,14),
		conv_std_logic_vector(3405,14),
		conv_std_logic_vector(3399,14),
		conv_std_logic_vector(3394,14),
		conv_std_logic_vector(3388,14),
		conv_std_logic_vector(3382,14),
		conv_std_logic_vector(3377,14),
		conv_std_logic_vector(3371,14),
		conv_std_logic_vector(3365,14),
		conv_std_logic_vector(3359,14),
		conv_std_logic_vector(3354,14),
		conv_std_logic_vector(3348,14),
		conv_std_logic_vector(3342,14),
		conv_std_logic_vector(3336,14),
		conv_std_logic_vector(3331,14),
		conv_std_logic_vector(3325,14),
		conv_std_logic_vector(3319,14),
		conv_std_logic_vector(3313,14),
		conv_std_logic_vector(3308,14),
		conv_std_logic_vector(3302,14),
		conv_std_logic_vector(3296,14),
		conv_std_logic_vector(3290,14),
		conv_std_logic_vector(3285,14),
		conv_std_logic_vector(3279,14),
		conv_std_logic_vector(3273,14),
		conv_std_logic_vector(3267,14),
		conv_std_logic_vector(3262,14),
		conv_std_logic_vector(3256,14),
		conv_std_logic_vector(3250,14),
		conv_std_logic_vector(3244,14),
		conv_std_logic_vector(3239,14),
		conv_std_logic_vector(3233,14),
		conv_std_logic_vector(3227,14),
		conv_std_logic_vector(3221,14),
		conv_std_logic_vector(3216,14),
		conv_std_logic_vector(3210,14),
		conv_std_logic_vector(3204,14),
		conv_std_logic_vector(3198,14),
		conv_std_logic_vector(3192,14),
		conv_std_logic_vector(3187,14),
		conv_std_logic_vector(3181,14),
		conv_std_logic_vector(3175,14),
		conv_std_logic_vector(3169,14),
		conv_std_logic_vector(3163,14),
		conv_std_logic_vector(3158,14),
		conv_std_logic_vector(3152,14),
		conv_std_logic_vector(3146,14),
		conv_std_logic_vector(3140,14),
		conv_std_logic_vector(3134,14),
		conv_std_logic_vector(3129,14),
		conv_std_logic_vector(3123,14),
		conv_std_logic_vector(3117,14),
		conv_std_logic_vector(3111,14),
		conv_std_logic_vector(3105,14),
		conv_std_logic_vector(3100,14),
		conv_std_logic_vector(3094,14),
		conv_std_logic_vector(3088,14),
		conv_std_logic_vector(3082,14),
		conv_std_logic_vector(3076,14),
		conv_std_logic_vector(3070,14),
		conv_std_logic_vector(3065,14),
		conv_std_logic_vector(3059,14),
		conv_std_logic_vector(3053,14),
		conv_std_logic_vector(3047,14),
		conv_std_logic_vector(3041,14),
		conv_std_logic_vector(3035,14),
		conv_std_logic_vector(3030,14),
		conv_std_logic_vector(3024,14),
		conv_std_logic_vector(3018,14),
		conv_std_logic_vector(3012,14),
		conv_std_logic_vector(3006,14),
		conv_std_logic_vector(3000,14),
		conv_std_logic_vector(2995,14),
		conv_std_logic_vector(2989,14),
		conv_std_logic_vector(2983,14),
		conv_std_logic_vector(2977,14),
		conv_std_logic_vector(2971,14),
		conv_std_logic_vector(2965,14),
		conv_std_logic_vector(2959,14),
		conv_std_logic_vector(2954,14),
		conv_std_logic_vector(2948,14),
		conv_std_logic_vector(2942,14),
		conv_std_logic_vector(2936,14),
		conv_std_logic_vector(2930,14),
		conv_std_logic_vector(2924,14),
		conv_std_logic_vector(2918,14),
		conv_std_logic_vector(2913,14),
		conv_std_logic_vector(2907,14),
		conv_std_logic_vector(2901,14),
		conv_std_logic_vector(2895,14),
		conv_std_logic_vector(2889,14),
		conv_std_logic_vector(2883,14),
		conv_std_logic_vector(2877,14),
		conv_std_logic_vector(2871,14),
		conv_std_logic_vector(2866,14),
		conv_std_logic_vector(2860,14),
		conv_std_logic_vector(2854,14),
		conv_std_logic_vector(2848,14),
		conv_std_logic_vector(2842,14),
		conv_std_logic_vector(2836,14),
		conv_std_logic_vector(2830,14),
		conv_std_logic_vector(2824,14),
		conv_std_logic_vector(2818,14),
		conv_std_logic_vector(2812,14),
		conv_std_logic_vector(2807,14),
		conv_std_logic_vector(2801,14),
		conv_std_logic_vector(2795,14),
		conv_std_logic_vector(2789,14),
		conv_std_logic_vector(2783,14),
		conv_std_logic_vector(2777,14),
		conv_std_logic_vector(2771,14),
		conv_std_logic_vector(2765,14),
		conv_std_logic_vector(2759,14),
		conv_std_logic_vector(2753,14),
		conv_std_logic_vector(2747,14),
		conv_std_logic_vector(2742,14),
		conv_std_logic_vector(2736,14),
		conv_std_logic_vector(2730,14),
		conv_std_logic_vector(2724,14),
		conv_std_logic_vector(2718,14),
		conv_std_logic_vector(2712,14),
		conv_std_logic_vector(2706,14),
		conv_std_logic_vector(2700,14),
		conv_std_logic_vector(2694,14),
		conv_std_logic_vector(2688,14),
		conv_std_logic_vector(2682,14),
		conv_std_logic_vector(2676,14),
		conv_std_logic_vector(2670,14),
		conv_std_logic_vector(2664,14),
		conv_std_logic_vector(2658,14),
		conv_std_logic_vector(2653,14),
		conv_std_logic_vector(2647,14),
		conv_std_logic_vector(2641,14),
		conv_std_logic_vector(2635,14),
		conv_std_logic_vector(2629,14),
		conv_std_logic_vector(2623,14),
		conv_std_logic_vector(2617,14),
		conv_std_logic_vector(2611,14),
		conv_std_logic_vector(2605,14),
		conv_std_logic_vector(2599,14),
		conv_std_logic_vector(2593,14),
		conv_std_logic_vector(2587,14),
		conv_std_logic_vector(2581,14),
		conv_std_logic_vector(2575,14),
		conv_std_logic_vector(2569,14),
		conv_std_logic_vector(2563,14),
		conv_std_logic_vector(2557,14),
		conv_std_logic_vector(2551,14),
		conv_std_logic_vector(2545,14),
		conv_std_logic_vector(2539,14),
		conv_std_logic_vector(2533,14),
		conv_std_logic_vector(2527,14),
		conv_std_logic_vector(2521,14),
		conv_std_logic_vector(2515,14),
		conv_std_logic_vector(2509,14),
		conv_std_logic_vector(2503,14),
		conv_std_logic_vector(2497,14),
		conv_std_logic_vector(2491,14),
		conv_std_logic_vector(2486,14),
		conv_std_logic_vector(2480,14),
		conv_std_logic_vector(2474,14),
		conv_std_logic_vector(2468,14),
		conv_std_logic_vector(2462,14),
		conv_std_logic_vector(2456,14),
		conv_std_logic_vector(2450,14),
		conv_std_logic_vector(2444,14),
		conv_std_logic_vector(2438,14),
		conv_std_logic_vector(2432,14),
		conv_std_logic_vector(2426,14),
		conv_std_logic_vector(2420,14),
		conv_std_logic_vector(2414,14),
		conv_std_logic_vector(2408,14),
		conv_std_logic_vector(2402,14),
		conv_std_logic_vector(2396,14),
		conv_std_logic_vector(2390,14),
		conv_std_logic_vector(2384,14),
		conv_std_logic_vector(2378,14),
		conv_std_logic_vector(2371,14),
		conv_std_logic_vector(2365,14),
		conv_std_logic_vector(2359,14),
		conv_std_logic_vector(2353,14),
		conv_std_logic_vector(2347,14),
		conv_std_logic_vector(2341,14),
		conv_std_logic_vector(2335,14),
		conv_std_logic_vector(2329,14),
		conv_std_logic_vector(2323,14),
		conv_std_logic_vector(2317,14),
		conv_std_logic_vector(2311,14),
		conv_std_logic_vector(2305,14),
		conv_std_logic_vector(2299,14),
		conv_std_logic_vector(2293,14),
		conv_std_logic_vector(2287,14),
		conv_std_logic_vector(2281,14),
		conv_std_logic_vector(2275,14),
		conv_std_logic_vector(2269,14),
		conv_std_logic_vector(2263,14),
		conv_std_logic_vector(2257,14),
		conv_std_logic_vector(2251,14),
		conv_std_logic_vector(2245,14),
		conv_std_logic_vector(2239,14),
		conv_std_logic_vector(2233,14),
		conv_std_logic_vector(2227,14),
		conv_std_logic_vector(2221,14),
		conv_std_logic_vector(2215,14),
		conv_std_logic_vector(2209,14),
		conv_std_logic_vector(2203,14),
		conv_std_logic_vector(2197,14),
		conv_std_logic_vector(2190,14),
		conv_std_logic_vector(2184,14),
		conv_std_logic_vector(2178,14),
		conv_std_logic_vector(2172,14),
		conv_std_logic_vector(2166,14),
		conv_std_logic_vector(2160,14),
		conv_std_logic_vector(2154,14),
		conv_std_logic_vector(2148,14),
		conv_std_logic_vector(2142,14),
		conv_std_logic_vector(2136,14),
		conv_std_logic_vector(2130,14),
		conv_std_logic_vector(2124,14),
		conv_std_logic_vector(2118,14),
		conv_std_logic_vector(2112,14),
		conv_std_logic_vector(2106,14),
		conv_std_logic_vector(2100,14),
		conv_std_logic_vector(2093,14),
		conv_std_logic_vector(2087,14),
		conv_std_logic_vector(2081,14),
		conv_std_logic_vector(2075,14),
		conv_std_logic_vector(2069,14),
		conv_std_logic_vector(2063,14),
		conv_std_logic_vector(2057,14),
		conv_std_logic_vector(2051,14),
		conv_std_logic_vector(2045,14),
		conv_std_logic_vector(2039,14),
		conv_std_logic_vector(2033,14),
		conv_std_logic_vector(2027,14),
		conv_std_logic_vector(2020,14),
		conv_std_logic_vector(2014,14),
		conv_std_logic_vector(2008,14),
		conv_std_logic_vector(2002,14),
		conv_std_logic_vector(1996,14),
		conv_std_logic_vector(1990,14),
		conv_std_logic_vector(1984,14),
		conv_std_logic_vector(1978,14),
		conv_std_logic_vector(1972,14),
		conv_std_logic_vector(1966,14),
		conv_std_logic_vector(1960,14),
		conv_std_logic_vector(1953,14),
		conv_std_logic_vector(1947,14),
		conv_std_logic_vector(1941,14),
		conv_std_logic_vector(1935,14),
		conv_std_logic_vector(1929,14),
		conv_std_logic_vector(1923,14),
		conv_std_logic_vector(1917,14),
		conv_std_logic_vector(1911,14),
		conv_std_logic_vector(1905,14),
		conv_std_logic_vector(1898,14),
		conv_std_logic_vector(1892,14),
		conv_std_logic_vector(1886,14),
		conv_std_logic_vector(1880,14),
		conv_std_logic_vector(1874,14),
		conv_std_logic_vector(1868,14),
		conv_std_logic_vector(1862,14),
		conv_std_logic_vector(1856,14),
		conv_std_logic_vector(1850,14),
		conv_std_logic_vector(1843,14),
		conv_std_logic_vector(1837,14),
		conv_std_logic_vector(1831,14),
		conv_std_logic_vector(1825,14),
		conv_std_logic_vector(1819,14),
		conv_std_logic_vector(1813,14),
		conv_std_logic_vector(1807,14),
		conv_std_logic_vector(1801,14),
		conv_std_logic_vector(1794,14),
		conv_std_logic_vector(1788,14),
		conv_std_logic_vector(1782,14),
		conv_std_logic_vector(1776,14),
		conv_std_logic_vector(1770,14),
		conv_std_logic_vector(1764,14),
		conv_std_logic_vector(1758,14),
		conv_std_logic_vector(1751,14),
		conv_std_logic_vector(1745,14),
		conv_std_logic_vector(1739,14),
		conv_std_logic_vector(1733,14),
		conv_std_logic_vector(1727,14),
		conv_std_logic_vector(1721,14),
		conv_std_logic_vector(1715,14),
		conv_std_logic_vector(1708,14),
		conv_std_logic_vector(1702,14),
		conv_std_logic_vector(1696,14),
		conv_std_logic_vector(1690,14),
		conv_std_logic_vector(1684,14),
		conv_std_logic_vector(1678,14),
		conv_std_logic_vector(1672,14),
		conv_std_logic_vector(1665,14),
		conv_std_logic_vector(1659,14),
		conv_std_logic_vector(1653,14),
		conv_std_logic_vector(1647,14),
		conv_std_logic_vector(1641,14),
		conv_std_logic_vector(1635,14),
		conv_std_logic_vector(1628,14),
		conv_std_logic_vector(1622,14),
		conv_std_logic_vector(1616,14),
		conv_std_logic_vector(1610,14),
		conv_std_logic_vector(1604,14),
		conv_std_logic_vector(1598,14),
		conv_std_logic_vector(1592,14),
		conv_std_logic_vector(1585,14),
		conv_std_logic_vector(1579,14),
		conv_std_logic_vector(1573,14),
		conv_std_logic_vector(1567,14),
		conv_std_logic_vector(1561,14),
		conv_std_logic_vector(1555,14),
		conv_std_logic_vector(1548,14),
		conv_std_logic_vector(1542,14),
		conv_std_logic_vector(1536,14),
		conv_std_logic_vector(1530,14),
		conv_std_logic_vector(1524,14),
		conv_std_logic_vector(1517,14),
		conv_std_logic_vector(1511,14),
		conv_std_logic_vector(1505,14),
		conv_std_logic_vector(1499,14),
		conv_std_logic_vector(1493,14),
		conv_std_logic_vector(1487,14),
		conv_std_logic_vector(1480,14),
		conv_std_logic_vector(1474,14),
		conv_std_logic_vector(1468,14),
		conv_std_logic_vector(1462,14),
		conv_std_logic_vector(1456,14),
		conv_std_logic_vector(1450,14),
		conv_std_logic_vector(1443,14),
		conv_std_logic_vector(1437,14),
		conv_std_logic_vector(1431,14),
		conv_std_logic_vector(1425,14),
		conv_std_logic_vector(1419,14),
		conv_std_logic_vector(1412,14),
		conv_std_logic_vector(1406,14),
		conv_std_logic_vector(1400,14),
		conv_std_logic_vector(1394,14),
		conv_std_logic_vector(1388,14),
		conv_std_logic_vector(1381,14),
		conv_std_logic_vector(1375,14),
		conv_std_logic_vector(1369,14),
		conv_std_logic_vector(1363,14),
		conv_std_logic_vector(1357,14),
		conv_std_logic_vector(1350,14),
		conv_std_logic_vector(1344,14),
		conv_std_logic_vector(1338,14),
		conv_std_logic_vector(1332,14),
		conv_std_logic_vector(1326,14),
		conv_std_logic_vector(1319,14),
		conv_std_logic_vector(1313,14),
		conv_std_logic_vector(1307,14),
		conv_std_logic_vector(1301,14),
		conv_std_logic_vector(1295,14),
		conv_std_logic_vector(1288,14),
		conv_std_logic_vector(1282,14),
		conv_std_logic_vector(1276,14),
		conv_std_logic_vector(1270,14),
		conv_std_logic_vector(1264,14),
		conv_std_logic_vector(1257,14),
		conv_std_logic_vector(1251,14),
		conv_std_logic_vector(1245,14),
		conv_std_logic_vector(1239,14),
		conv_std_logic_vector(1233,14),
		conv_std_logic_vector(1226,14),
		conv_std_logic_vector(1220,14),
		conv_std_logic_vector(1214,14),
		conv_std_logic_vector(1208,14),
		conv_std_logic_vector(1202,14),
		conv_std_logic_vector(1195,14),
		conv_std_logic_vector(1189,14),
		conv_std_logic_vector(1183,14),
		conv_std_logic_vector(1177,14),
		conv_std_logic_vector(1170,14),
		conv_std_logic_vector(1164,14),
		conv_std_logic_vector(1158,14),
		conv_std_logic_vector(1152,14),
		conv_std_logic_vector(1146,14),
		conv_std_logic_vector(1139,14),
		conv_std_logic_vector(1133,14),
		conv_std_logic_vector(1127,14),
		conv_std_logic_vector(1121,14),
		conv_std_logic_vector(1114,14),
		conv_std_logic_vector(1108,14),
		conv_std_logic_vector(1102,14),
		conv_std_logic_vector(1096,14),
		conv_std_logic_vector(1090,14),
		conv_std_logic_vector(1083,14),
		conv_std_logic_vector(1077,14),
		conv_std_logic_vector(1071,14),
		conv_std_logic_vector(1065,14),
		conv_std_logic_vector(1058,14),
		conv_std_logic_vector(1052,14),
		conv_std_logic_vector(1046,14),
		conv_std_logic_vector(1040,14),
		conv_std_logic_vector(1033,14),
		conv_std_logic_vector(1027,14),
		conv_std_logic_vector(1021,14),
		conv_std_logic_vector(1015,14),
		conv_std_logic_vector(1009,14),
		conv_std_logic_vector(1002,14),
		conv_std_logic_vector(996,14),
		conv_std_logic_vector(990,14),
		conv_std_logic_vector(984,14),
		conv_std_logic_vector(977,14),
		conv_std_logic_vector(971,14),
		conv_std_logic_vector(965,14),
		conv_std_logic_vector(959,14),
		conv_std_logic_vector(952,14),
		conv_std_logic_vector(946,14),
		conv_std_logic_vector(940,14),
		conv_std_logic_vector(934,14),
		conv_std_logic_vector(927,14),
		conv_std_logic_vector(921,14),
		conv_std_logic_vector(915,14),
		conv_std_logic_vector(909,14),
		conv_std_logic_vector(902,14),
		conv_std_logic_vector(896,14),
		conv_std_logic_vector(890,14),
		conv_std_logic_vector(884,14),
		conv_std_logic_vector(877,14),
		conv_std_logic_vector(871,14),
		conv_std_logic_vector(865,14),
		conv_std_logic_vector(859,14),
		conv_std_logic_vector(852,14),
		conv_std_logic_vector(846,14),
		conv_std_logic_vector(840,14),
		conv_std_logic_vector(834,14),
		conv_std_logic_vector(827,14),
		conv_std_logic_vector(821,14),
		conv_std_logic_vector(815,14),
		conv_std_logic_vector(809,14),
		conv_std_logic_vector(802,14),
		conv_std_logic_vector(796,14),
		conv_std_logic_vector(790,14),
		conv_std_logic_vector(784,14),
		conv_std_logic_vector(777,14),
		conv_std_logic_vector(771,14),
		conv_std_logic_vector(765,14),
		conv_std_logic_vector(759,14),
		conv_std_logic_vector(752,14),
		conv_std_logic_vector(746,14),
		conv_std_logic_vector(740,14),
		conv_std_logic_vector(734,14),
		conv_std_logic_vector(727,14),
		conv_std_logic_vector(721,14),
		conv_std_logic_vector(715,14),
		conv_std_logic_vector(709,14),
		conv_std_logic_vector(702,14),
		conv_std_logic_vector(696,14),
		conv_std_logic_vector(690,14),
		conv_std_logic_vector(684,14),
		conv_std_logic_vector(677,14),
		conv_std_logic_vector(671,14),
		conv_std_logic_vector(665,14),
		conv_std_logic_vector(659,14),
		conv_std_logic_vector(652,14),
		conv_std_logic_vector(646,14),
		conv_std_logic_vector(640,14),
		conv_std_logic_vector(633,14),
		conv_std_logic_vector(627,14),
		conv_std_logic_vector(621,14),
		conv_std_logic_vector(615,14),
		conv_std_logic_vector(608,14),
		conv_std_logic_vector(602,14),
		conv_std_logic_vector(596,14),
		conv_std_logic_vector(590,14),
		conv_std_logic_vector(583,14),
		conv_std_logic_vector(577,14),
		conv_std_logic_vector(571,14),
		conv_std_logic_vector(565,14),
		conv_std_logic_vector(558,14),
		conv_std_logic_vector(552,14),
		conv_std_logic_vector(546,14),
		conv_std_logic_vector(539,14),
		conv_std_logic_vector(533,14),
		conv_std_logic_vector(527,14),
		conv_std_logic_vector(521,14),
		conv_std_logic_vector(514,14),
		conv_std_logic_vector(508,14),
		conv_std_logic_vector(502,14),
		conv_std_logic_vector(496,14),
		conv_std_logic_vector(489,14),
		conv_std_logic_vector(483,14),
		conv_std_logic_vector(477,14),
		conv_std_logic_vector(470,14),
		conv_std_logic_vector(464,14),
		conv_std_logic_vector(458,14),
		conv_std_logic_vector(452,14),
		conv_std_logic_vector(445,14),
		conv_std_logic_vector(439,14),
		conv_std_logic_vector(433,14),
		conv_std_logic_vector(427,14),
		conv_std_logic_vector(420,14),
		conv_std_logic_vector(414,14),
		conv_std_logic_vector(408,14),
		conv_std_logic_vector(401,14),
		conv_std_logic_vector(395,14),
		conv_std_logic_vector(389,14),
		conv_std_logic_vector(383,14),
		conv_std_logic_vector(376,14),
		conv_std_logic_vector(370,14),
		conv_std_logic_vector(364,14),
		conv_std_logic_vector(358,14),
		conv_std_logic_vector(351,14),
		conv_std_logic_vector(345,14),
		conv_std_logic_vector(339,14),
		conv_std_logic_vector(332,14),
		conv_std_logic_vector(326,14),
		conv_std_logic_vector(320,14),
		conv_std_logic_vector(314,14),
		conv_std_logic_vector(307,14),
		conv_std_logic_vector(301,14),
		conv_std_logic_vector(295,14),
		conv_std_logic_vector(288,14),
		conv_std_logic_vector(282,14),
		conv_std_logic_vector(276,14),
		conv_std_logic_vector(270,14),
		conv_std_logic_vector(263,14),
		conv_std_logic_vector(257,14),
		conv_std_logic_vector(251,14),
		conv_std_logic_vector(245,14),
		conv_std_logic_vector(238,14),
		conv_std_logic_vector(232,14),
		conv_std_logic_vector(226,14),
		conv_std_logic_vector(219,14),
		conv_std_logic_vector(213,14),
		conv_std_logic_vector(207,14),
		conv_std_logic_vector(201,14),
		conv_std_logic_vector(194,14),
		conv_std_logic_vector(188,14),
		conv_std_logic_vector(182,14),
		conv_std_logic_vector(175,14),
		conv_std_logic_vector(169,14),
		conv_std_logic_vector(163,14),
		conv_std_logic_vector(157,14),
		conv_std_logic_vector(150,14),
		conv_std_logic_vector(144,14),
		conv_std_logic_vector(138,14),
		conv_std_logic_vector(131,14),
		conv_std_logic_vector(125,14),
		conv_std_logic_vector(119,14),
		conv_std_logic_vector(113,14),
		conv_std_logic_vector(106,14),
		conv_std_logic_vector(100,14),
		conv_std_logic_vector(94,14),
		conv_std_logic_vector(87,14),
		conv_std_logic_vector(81,14),
		conv_std_logic_vector(75,14),
		conv_std_logic_vector(69,14),
		conv_std_logic_vector(62,14),
		conv_std_logic_vector(56,14),
		conv_std_logic_vector(50,14),
		conv_std_logic_vector(43,14),
		conv_std_logic_vector(37,14),
		conv_std_logic_vector(31,14),
		conv_std_logic_vector(25,14),
		conv_std_logic_vector(18,14),
		conv_std_logic_vector(12,14),
		conv_std_logic_vector(6,14),
		conv_std_logic_vector(0,14),
		conv_std_logic_vector(-6,14),
		conv_std_logic_vector(-12,14),
		conv_std_logic_vector(-18,14),
		conv_std_logic_vector(-25,14),
		conv_std_logic_vector(-31,14),
		conv_std_logic_vector(-37,14),
		conv_std_logic_vector(-43,14),
		conv_std_logic_vector(-50,14),
		conv_std_logic_vector(-56,14),
		conv_std_logic_vector(-62,14),
		conv_std_logic_vector(-69,14),
		conv_std_logic_vector(-75,14),
		conv_std_logic_vector(-81,14),
		conv_std_logic_vector(-87,14),
		conv_std_logic_vector(-94,14),
		conv_std_logic_vector(-100,14),
		conv_std_logic_vector(-106,14),
		conv_std_logic_vector(-113,14),
		conv_std_logic_vector(-119,14),
		conv_std_logic_vector(-125,14),
		conv_std_logic_vector(-131,14),
		conv_std_logic_vector(-138,14),
		conv_std_logic_vector(-144,14),
		conv_std_logic_vector(-150,14),
		conv_std_logic_vector(-157,14),
		conv_std_logic_vector(-163,14),
		conv_std_logic_vector(-169,14),
		conv_std_logic_vector(-175,14),
		conv_std_logic_vector(-182,14),
		conv_std_logic_vector(-188,14),
		conv_std_logic_vector(-194,14),
		conv_std_logic_vector(-201,14),
		conv_std_logic_vector(-207,14),
		conv_std_logic_vector(-213,14),
		conv_std_logic_vector(-219,14),
		conv_std_logic_vector(-226,14),
		conv_std_logic_vector(-232,14),
		conv_std_logic_vector(-238,14),
		conv_std_logic_vector(-245,14),
		conv_std_logic_vector(-251,14),
		conv_std_logic_vector(-257,14),
		conv_std_logic_vector(-263,14),
		conv_std_logic_vector(-270,14),
		conv_std_logic_vector(-276,14),
		conv_std_logic_vector(-282,14),
		conv_std_logic_vector(-288,14),
		conv_std_logic_vector(-295,14),
		conv_std_logic_vector(-301,14),
		conv_std_logic_vector(-307,14),
		conv_std_logic_vector(-314,14),
		conv_std_logic_vector(-320,14),
		conv_std_logic_vector(-326,14),
		conv_std_logic_vector(-332,14),
		conv_std_logic_vector(-339,14),
		conv_std_logic_vector(-345,14),
		conv_std_logic_vector(-351,14),
		conv_std_logic_vector(-358,14),
		conv_std_logic_vector(-364,14),
		conv_std_logic_vector(-370,14),
		conv_std_logic_vector(-376,14),
		conv_std_logic_vector(-383,14),
		conv_std_logic_vector(-389,14),
		conv_std_logic_vector(-395,14),
		conv_std_logic_vector(-401,14),
		conv_std_logic_vector(-408,14),
		conv_std_logic_vector(-414,14),
		conv_std_logic_vector(-420,14),
		conv_std_logic_vector(-427,14),
		conv_std_logic_vector(-433,14),
		conv_std_logic_vector(-439,14),
		conv_std_logic_vector(-445,14),
		conv_std_logic_vector(-452,14),
		conv_std_logic_vector(-458,14),
		conv_std_logic_vector(-464,14),
		conv_std_logic_vector(-470,14),
		conv_std_logic_vector(-477,14),
		conv_std_logic_vector(-483,14),
		conv_std_logic_vector(-489,14),
		conv_std_logic_vector(-496,14),
		conv_std_logic_vector(-502,14),
		conv_std_logic_vector(-508,14),
		conv_std_logic_vector(-514,14),
		conv_std_logic_vector(-521,14),
		conv_std_logic_vector(-527,14),
		conv_std_logic_vector(-533,14),
		conv_std_logic_vector(-539,14),
		conv_std_logic_vector(-546,14),
		conv_std_logic_vector(-552,14),
		conv_std_logic_vector(-558,14),
		conv_std_logic_vector(-565,14),
		conv_std_logic_vector(-571,14),
		conv_std_logic_vector(-577,14),
		conv_std_logic_vector(-583,14),
		conv_std_logic_vector(-590,14),
		conv_std_logic_vector(-596,14),
		conv_std_logic_vector(-602,14),
		conv_std_logic_vector(-608,14),
		conv_std_logic_vector(-615,14),
		conv_std_logic_vector(-621,14),
		conv_std_logic_vector(-627,14),
		conv_std_logic_vector(-633,14),
		conv_std_logic_vector(-640,14),
		conv_std_logic_vector(-646,14),
		conv_std_logic_vector(-652,14),
		conv_std_logic_vector(-659,14),
		conv_std_logic_vector(-665,14),
		conv_std_logic_vector(-671,14),
		conv_std_logic_vector(-677,14),
		conv_std_logic_vector(-684,14),
		conv_std_logic_vector(-690,14),
		conv_std_logic_vector(-696,14),
		conv_std_logic_vector(-702,14),
		conv_std_logic_vector(-709,14),
		conv_std_logic_vector(-715,14),
		conv_std_logic_vector(-721,14),
		conv_std_logic_vector(-727,14),
		conv_std_logic_vector(-734,14),
		conv_std_logic_vector(-740,14),
		conv_std_logic_vector(-746,14),
		conv_std_logic_vector(-752,14),
		conv_std_logic_vector(-759,14),
		conv_std_logic_vector(-765,14),
		conv_std_logic_vector(-771,14),
		conv_std_logic_vector(-777,14),
		conv_std_logic_vector(-784,14),
		conv_std_logic_vector(-790,14),
		conv_std_logic_vector(-796,14),
		conv_std_logic_vector(-802,14),
		conv_std_logic_vector(-809,14),
		conv_std_logic_vector(-815,14),
		conv_std_logic_vector(-821,14),
		conv_std_logic_vector(-827,14),
		conv_std_logic_vector(-834,14),
		conv_std_logic_vector(-840,14),
		conv_std_logic_vector(-846,14),
		conv_std_logic_vector(-852,14),
		conv_std_logic_vector(-859,14),
		conv_std_logic_vector(-865,14),
		conv_std_logic_vector(-871,14),
		conv_std_logic_vector(-877,14),
		conv_std_logic_vector(-884,14),
		conv_std_logic_vector(-890,14),
		conv_std_logic_vector(-896,14),
		conv_std_logic_vector(-902,14),
		conv_std_logic_vector(-909,14),
		conv_std_logic_vector(-915,14),
		conv_std_logic_vector(-921,14),
		conv_std_logic_vector(-927,14),
		conv_std_logic_vector(-934,14),
		conv_std_logic_vector(-940,14),
		conv_std_logic_vector(-946,14),
		conv_std_logic_vector(-952,14),
		conv_std_logic_vector(-959,14),
		conv_std_logic_vector(-965,14),
		conv_std_logic_vector(-971,14),
		conv_std_logic_vector(-977,14),
		conv_std_logic_vector(-984,14),
		conv_std_logic_vector(-990,14),
		conv_std_logic_vector(-996,14),
		conv_std_logic_vector(-1002,14),
		conv_std_logic_vector(-1009,14),
		conv_std_logic_vector(-1015,14),
		conv_std_logic_vector(-1021,14),
		conv_std_logic_vector(-1027,14),
		conv_std_logic_vector(-1033,14),
		conv_std_logic_vector(-1040,14),
		conv_std_logic_vector(-1046,14),
		conv_std_logic_vector(-1052,14),
		conv_std_logic_vector(-1058,14),
		conv_std_logic_vector(-1065,14),
		conv_std_logic_vector(-1071,14),
		conv_std_logic_vector(-1077,14),
		conv_std_logic_vector(-1083,14),
		conv_std_logic_vector(-1090,14),
		conv_std_logic_vector(-1096,14),
		conv_std_logic_vector(-1102,14),
		conv_std_logic_vector(-1108,14),
		conv_std_logic_vector(-1114,14),
		conv_std_logic_vector(-1121,14),
		conv_std_logic_vector(-1127,14),
		conv_std_logic_vector(-1133,14),
		conv_std_logic_vector(-1139,14),
		conv_std_logic_vector(-1146,14),
		conv_std_logic_vector(-1152,14),
		conv_std_logic_vector(-1158,14),
		conv_std_logic_vector(-1164,14),
		conv_std_logic_vector(-1170,14),
		conv_std_logic_vector(-1177,14),
		conv_std_logic_vector(-1183,14),
		conv_std_logic_vector(-1189,14),
		conv_std_logic_vector(-1195,14),
		conv_std_logic_vector(-1202,14),
		conv_std_logic_vector(-1208,14),
		conv_std_logic_vector(-1214,14),
		conv_std_logic_vector(-1220,14),
		conv_std_logic_vector(-1226,14),
		conv_std_logic_vector(-1233,14),
		conv_std_logic_vector(-1239,14),
		conv_std_logic_vector(-1245,14),
		conv_std_logic_vector(-1251,14),
		conv_std_logic_vector(-1257,14),
		conv_std_logic_vector(-1264,14),
		conv_std_logic_vector(-1270,14),
		conv_std_logic_vector(-1276,14),
		conv_std_logic_vector(-1282,14),
		conv_std_logic_vector(-1288,14),
		conv_std_logic_vector(-1295,14),
		conv_std_logic_vector(-1301,14),
		conv_std_logic_vector(-1307,14),
		conv_std_logic_vector(-1313,14),
		conv_std_logic_vector(-1319,14),
		conv_std_logic_vector(-1326,14),
		conv_std_logic_vector(-1332,14),
		conv_std_logic_vector(-1338,14),
		conv_std_logic_vector(-1344,14),
		conv_std_logic_vector(-1350,14),
		conv_std_logic_vector(-1357,14),
		conv_std_logic_vector(-1363,14),
		conv_std_logic_vector(-1369,14),
		conv_std_logic_vector(-1375,14),
		conv_std_logic_vector(-1381,14),
		conv_std_logic_vector(-1388,14),
		conv_std_logic_vector(-1394,14),
		conv_std_logic_vector(-1400,14),
		conv_std_logic_vector(-1406,14),
		conv_std_logic_vector(-1412,14),
		conv_std_logic_vector(-1419,14),
		conv_std_logic_vector(-1425,14),
		conv_std_logic_vector(-1431,14),
		conv_std_logic_vector(-1437,14),
		conv_std_logic_vector(-1443,14),
		conv_std_logic_vector(-1450,14),
		conv_std_logic_vector(-1456,14),
		conv_std_logic_vector(-1462,14),
		conv_std_logic_vector(-1468,14),
		conv_std_logic_vector(-1474,14),
		conv_std_logic_vector(-1480,14),
		conv_std_logic_vector(-1487,14),
		conv_std_logic_vector(-1493,14),
		conv_std_logic_vector(-1499,14),
		conv_std_logic_vector(-1505,14),
		conv_std_logic_vector(-1511,14),
		conv_std_logic_vector(-1517,14),
		conv_std_logic_vector(-1524,14),
		conv_std_logic_vector(-1530,14),
		conv_std_logic_vector(-1536,14),
		conv_std_logic_vector(-1542,14),
		conv_std_logic_vector(-1548,14),
		conv_std_logic_vector(-1555,14),
		conv_std_logic_vector(-1561,14),
		conv_std_logic_vector(-1567,14),
		conv_std_logic_vector(-1573,14),
		conv_std_logic_vector(-1579,14),
		conv_std_logic_vector(-1585,14),
		conv_std_logic_vector(-1592,14),
		conv_std_logic_vector(-1598,14),
		conv_std_logic_vector(-1604,14),
		conv_std_logic_vector(-1610,14),
		conv_std_logic_vector(-1616,14),
		conv_std_logic_vector(-1622,14),
		conv_std_logic_vector(-1628,14),
		conv_std_logic_vector(-1635,14),
		conv_std_logic_vector(-1641,14),
		conv_std_logic_vector(-1647,14),
		conv_std_logic_vector(-1653,14),
		conv_std_logic_vector(-1659,14),
		conv_std_logic_vector(-1665,14),
		conv_std_logic_vector(-1672,14),
		conv_std_logic_vector(-1678,14),
		conv_std_logic_vector(-1684,14),
		conv_std_logic_vector(-1690,14),
		conv_std_logic_vector(-1696,14),
		conv_std_logic_vector(-1702,14),
		conv_std_logic_vector(-1708,14),
		conv_std_logic_vector(-1715,14),
		conv_std_logic_vector(-1721,14),
		conv_std_logic_vector(-1727,14),
		conv_std_logic_vector(-1733,14),
		conv_std_logic_vector(-1739,14),
		conv_std_logic_vector(-1745,14),
		conv_std_logic_vector(-1751,14),
		conv_std_logic_vector(-1758,14),
		conv_std_logic_vector(-1764,14),
		conv_std_logic_vector(-1770,14),
		conv_std_logic_vector(-1776,14),
		conv_std_logic_vector(-1782,14),
		conv_std_logic_vector(-1788,14),
		conv_std_logic_vector(-1794,14),
		conv_std_logic_vector(-1801,14),
		conv_std_logic_vector(-1807,14),
		conv_std_logic_vector(-1813,14),
		conv_std_logic_vector(-1819,14),
		conv_std_logic_vector(-1825,14),
		conv_std_logic_vector(-1831,14),
		conv_std_logic_vector(-1837,14),
		conv_std_logic_vector(-1843,14),
		conv_std_logic_vector(-1850,14),
		conv_std_logic_vector(-1856,14),
		conv_std_logic_vector(-1862,14),
		conv_std_logic_vector(-1868,14),
		conv_std_logic_vector(-1874,14),
		conv_std_logic_vector(-1880,14),
		conv_std_logic_vector(-1886,14),
		conv_std_logic_vector(-1892,14),
		conv_std_logic_vector(-1898,14),
		conv_std_logic_vector(-1905,14),
		conv_std_logic_vector(-1911,14),
		conv_std_logic_vector(-1917,14),
		conv_std_logic_vector(-1923,14),
		conv_std_logic_vector(-1929,14),
		conv_std_logic_vector(-1935,14),
		conv_std_logic_vector(-1941,14),
		conv_std_logic_vector(-1947,14),
		conv_std_logic_vector(-1953,14),
		conv_std_logic_vector(-1960,14),
		conv_std_logic_vector(-1966,14),
		conv_std_logic_vector(-1972,14),
		conv_std_logic_vector(-1978,14),
		conv_std_logic_vector(-1984,14),
		conv_std_logic_vector(-1990,14),
		conv_std_logic_vector(-1996,14),
		conv_std_logic_vector(-2002,14),
		conv_std_logic_vector(-2008,14),
		conv_std_logic_vector(-2014,14),
		conv_std_logic_vector(-2020,14),
		conv_std_logic_vector(-2027,14),
		conv_std_logic_vector(-2033,14),
		conv_std_logic_vector(-2039,14),
		conv_std_logic_vector(-2045,14),
		conv_std_logic_vector(-2051,14),
		conv_std_logic_vector(-2057,14),
		conv_std_logic_vector(-2063,14),
		conv_std_logic_vector(-2069,14),
		conv_std_logic_vector(-2075,14),
		conv_std_logic_vector(-2081,14),
		conv_std_logic_vector(-2087,14),
		conv_std_logic_vector(-2093,14),
		conv_std_logic_vector(-2100,14),
		conv_std_logic_vector(-2106,14),
		conv_std_logic_vector(-2112,14),
		conv_std_logic_vector(-2118,14),
		conv_std_logic_vector(-2124,14),
		conv_std_logic_vector(-2130,14),
		conv_std_logic_vector(-2136,14),
		conv_std_logic_vector(-2142,14),
		conv_std_logic_vector(-2148,14),
		conv_std_logic_vector(-2154,14),
		conv_std_logic_vector(-2160,14),
		conv_std_logic_vector(-2166,14),
		conv_std_logic_vector(-2172,14),
		conv_std_logic_vector(-2178,14),
		conv_std_logic_vector(-2184,14),
		conv_std_logic_vector(-2190,14),
		conv_std_logic_vector(-2197,14),
		conv_std_logic_vector(-2203,14),
		conv_std_logic_vector(-2209,14),
		conv_std_logic_vector(-2215,14),
		conv_std_logic_vector(-2221,14),
		conv_std_logic_vector(-2227,14),
		conv_std_logic_vector(-2233,14),
		conv_std_logic_vector(-2239,14),
		conv_std_logic_vector(-2245,14),
		conv_std_logic_vector(-2251,14),
		conv_std_logic_vector(-2257,14),
		conv_std_logic_vector(-2263,14),
		conv_std_logic_vector(-2269,14),
		conv_std_logic_vector(-2275,14),
		conv_std_logic_vector(-2281,14),
		conv_std_logic_vector(-2287,14),
		conv_std_logic_vector(-2293,14),
		conv_std_logic_vector(-2299,14),
		conv_std_logic_vector(-2305,14),
		conv_std_logic_vector(-2311,14),
		conv_std_logic_vector(-2317,14),
		conv_std_logic_vector(-2323,14),
		conv_std_logic_vector(-2329,14),
		conv_std_logic_vector(-2335,14),
		conv_std_logic_vector(-2341,14),
		conv_std_logic_vector(-2347,14),
		conv_std_logic_vector(-2353,14),
		conv_std_logic_vector(-2359,14),
		conv_std_logic_vector(-2365,14),
		conv_std_logic_vector(-2371,14),
		conv_std_logic_vector(-2378,14),
		conv_std_logic_vector(-2384,14),
		conv_std_logic_vector(-2390,14),
		conv_std_logic_vector(-2396,14),
		conv_std_logic_vector(-2402,14),
		conv_std_logic_vector(-2408,14),
		conv_std_logic_vector(-2414,14),
		conv_std_logic_vector(-2420,14),
		conv_std_logic_vector(-2426,14),
		conv_std_logic_vector(-2432,14),
		conv_std_logic_vector(-2438,14),
		conv_std_logic_vector(-2444,14),
		conv_std_logic_vector(-2450,14),
		conv_std_logic_vector(-2456,14),
		conv_std_logic_vector(-2462,14),
		conv_std_logic_vector(-2468,14),
		conv_std_logic_vector(-2474,14),
		conv_std_logic_vector(-2480,14),
		conv_std_logic_vector(-2486,14),
		conv_std_logic_vector(-2491,14),
		conv_std_logic_vector(-2497,14),
		conv_std_logic_vector(-2503,14),
		conv_std_logic_vector(-2509,14),
		conv_std_logic_vector(-2515,14),
		conv_std_logic_vector(-2521,14),
		conv_std_logic_vector(-2527,14),
		conv_std_logic_vector(-2533,14),
		conv_std_logic_vector(-2539,14),
		conv_std_logic_vector(-2545,14),
		conv_std_logic_vector(-2551,14),
		conv_std_logic_vector(-2557,14),
		conv_std_logic_vector(-2563,14),
		conv_std_logic_vector(-2569,14),
		conv_std_logic_vector(-2575,14),
		conv_std_logic_vector(-2581,14),
		conv_std_logic_vector(-2587,14),
		conv_std_logic_vector(-2593,14),
		conv_std_logic_vector(-2599,14),
		conv_std_logic_vector(-2605,14),
		conv_std_logic_vector(-2611,14),
		conv_std_logic_vector(-2617,14),
		conv_std_logic_vector(-2623,14),
		conv_std_logic_vector(-2629,14),
		conv_std_logic_vector(-2635,14),
		conv_std_logic_vector(-2641,14),
		conv_std_logic_vector(-2647,14),
		conv_std_logic_vector(-2653,14),
		conv_std_logic_vector(-2658,14),
		conv_std_logic_vector(-2664,14),
		conv_std_logic_vector(-2670,14),
		conv_std_logic_vector(-2676,14),
		conv_std_logic_vector(-2682,14),
		conv_std_logic_vector(-2688,14),
		conv_std_logic_vector(-2694,14),
		conv_std_logic_vector(-2700,14),
		conv_std_logic_vector(-2706,14),
		conv_std_logic_vector(-2712,14),
		conv_std_logic_vector(-2718,14),
		conv_std_logic_vector(-2724,14),
		conv_std_logic_vector(-2730,14),
		conv_std_logic_vector(-2736,14),
		conv_std_logic_vector(-2742,14),
		conv_std_logic_vector(-2747,14),
		conv_std_logic_vector(-2753,14),
		conv_std_logic_vector(-2759,14),
		conv_std_logic_vector(-2765,14),
		conv_std_logic_vector(-2771,14),
		conv_std_logic_vector(-2777,14),
		conv_std_logic_vector(-2783,14),
		conv_std_logic_vector(-2789,14),
		conv_std_logic_vector(-2795,14),
		conv_std_logic_vector(-2801,14),
		conv_std_logic_vector(-2807,14),
		conv_std_logic_vector(-2812,14),
		conv_std_logic_vector(-2818,14),
		conv_std_logic_vector(-2824,14),
		conv_std_logic_vector(-2830,14),
		conv_std_logic_vector(-2836,14),
		conv_std_logic_vector(-2842,14),
		conv_std_logic_vector(-2848,14),
		conv_std_logic_vector(-2854,14),
		conv_std_logic_vector(-2860,14),
		conv_std_logic_vector(-2866,14),
		conv_std_logic_vector(-2871,14),
		conv_std_logic_vector(-2877,14),
		conv_std_logic_vector(-2883,14),
		conv_std_logic_vector(-2889,14),
		conv_std_logic_vector(-2895,14),
		conv_std_logic_vector(-2901,14),
		conv_std_logic_vector(-2907,14),
		conv_std_logic_vector(-2913,14),
		conv_std_logic_vector(-2918,14),
		conv_std_logic_vector(-2924,14),
		conv_std_logic_vector(-2930,14),
		conv_std_logic_vector(-2936,14),
		conv_std_logic_vector(-2942,14),
		conv_std_logic_vector(-2948,14),
		conv_std_logic_vector(-2954,14),
		conv_std_logic_vector(-2959,14),
		conv_std_logic_vector(-2965,14),
		conv_std_logic_vector(-2971,14),
		conv_std_logic_vector(-2977,14),
		conv_std_logic_vector(-2983,14),
		conv_std_logic_vector(-2989,14),
		conv_std_logic_vector(-2995,14),
		conv_std_logic_vector(-3000,14),
		conv_std_logic_vector(-3006,14),
		conv_std_logic_vector(-3012,14),
		conv_std_logic_vector(-3018,14),
		conv_std_logic_vector(-3024,14),
		conv_std_logic_vector(-3030,14),
		conv_std_logic_vector(-3035,14),
		conv_std_logic_vector(-3041,14),
		conv_std_logic_vector(-3047,14),
		conv_std_logic_vector(-3053,14),
		conv_std_logic_vector(-3059,14),
		conv_std_logic_vector(-3065,14),
		conv_std_logic_vector(-3070,14),
		conv_std_logic_vector(-3076,14),
		conv_std_logic_vector(-3082,14),
		conv_std_logic_vector(-3088,14),
		conv_std_logic_vector(-3094,14),
		conv_std_logic_vector(-3100,14),
		conv_std_logic_vector(-3105,14),
		conv_std_logic_vector(-3111,14),
		conv_std_logic_vector(-3117,14),
		conv_std_logic_vector(-3123,14),
		conv_std_logic_vector(-3129,14),
		conv_std_logic_vector(-3134,14),
		conv_std_logic_vector(-3140,14),
		conv_std_logic_vector(-3146,14),
		conv_std_logic_vector(-3152,14),
		conv_std_logic_vector(-3158,14),
		conv_std_logic_vector(-3163,14),
		conv_std_logic_vector(-3169,14),
		conv_std_logic_vector(-3175,14),
		conv_std_logic_vector(-3181,14),
		conv_std_logic_vector(-3187,14),
		conv_std_logic_vector(-3192,14),
		conv_std_logic_vector(-3198,14),
		conv_std_logic_vector(-3204,14),
		conv_std_logic_vector(-3210,14),
		conv_std_logic_vector(-3216,14),
		conv_std_logic_vector(-3221,14),
		conv_std_logic_vector(-3227,14),
		conv_std_logic_vector(-3233,14),
		conv_std_logic_vector(-3239,14),
		conv_std_logic_vector(-3244,14),
		conv_std_logic_vector(-3250,14),
		conv_std_logic_vector(-3256,14),
		conv_std_logic_vector(-3262,14),
		conv_std_logic_vector(-3267,14),
		conv_std_logic_vector(-3273,14),
		conv_std_logic_vector(-3279,14),
		conv_std_logic_vector(-3285,14),
		conv_std_logic_vector(-3290,14),
		conv_std_logic_vector(-3296,14),
		conv_std_logic_vector(-3302,14),
		conv_std_logic_vector(-3308,14),
		conv_std_logic_vector(-3313,14),
		conv_std_logic_vector(-3319,14),
		conv_std_logic_vector(-3325,14),
		conv_std_logic_vector(-3331,14),
		conv_std_logic_vector(-3336,14),
		conv_std_logic_vector(-3342,14),
		conv_std_logic_vector(-3348,14),
		conv_std_logic_vector(-3354,14),
		conv_std_logic_vector(-3359,14),
		conv_std_logic_vector(-3365,14),
		conv_std_logic_vector(-3371,14),
		conv_std_logic_vector(-3377,14),
		conv_std_logic_vector(-3382,14),
		conv_std_logic_vector(-3388,14),
		conv_std_logic_vector(-3394,14),
		conv_std_logic_vector(-3399,14),
		conv_std_logic_vector(-3405,14),
		conv_std_logic_vector(-3411,14),
		conv_std_logic_vector(-3417,14),
		conv_std_logic_vector(-3422,14),
		conv_std_logic_vector(-3428,14),
		conv_std_logic_vector(-3434,14),
		conv_std_logic_vector(-3439,14),
		conv_std_logic_vector(-3445,14),
		conv_std_logic_vector(-3451,14),
		conv_std_logic_vector(-3457,14),
		conv_std_logic_vector(-3462,14),
		conv_std_logic_vector(-3468,14),
		conv_std_logic_vector(-3474,14),
		conv_std_logic_vector(-3479,14),
		conv_std_logic_vector(-3485,14),
		conv_std_logic_vector(-3491,14),
		conv_std_logic_vector(-3496,14),
		conv_std_logic_vector(-3502,14),
		conv_std_logic_vector(-3508,14),
		conv_std_logic_vector(-3513,14),
		conv_std_logic_vector(-3519,14),
		conv_std_logic_vector(-3525,14),
		conv_std_logic_vector(-3530,14),
		conv_std_logic_vector(-3536,14),
		conv_std_logic_vector(-3542,14),
		conv_std_logic_vector(-3547,14),
		conv_std_logic_vector(-3553,14),
		conv_std_logic_vector(-3559,14),
		conv_std_logic_vector(-3564,14),
		conv_std_logic_vector(-3570,14),
		conv_std_logic_vector(-3576,14),
		conv_std_logic_vector(-3581,14),
		conv_std_logic_vector(-3587,14),
		conv_std_logic_vector(-3593,14),
		conv_std_logic_vector(-3598,14),
		conv_std_logic_vector(-3604,14),
		conv_std_logic_vector(-3610,14),
		conv_std_logic_vector(-3615,14),
		conv_std_logic_vector(-3621,14),
		conv_std_logic_vector(-3626,14),
		conv_std_logic_vector(-3632,14),
		conv_std_logic_vector(-3638,14),
		conv_std_logic_vector(-3643,14),
		conv_std_logic_vector(-3649,14),
		conv_std_logic_vector(-3655,14),
		conv_std_logic_vector(-3660,14),
		conv_std_logic_vector(-3666,14),
		conv_std_logic_vector(-3671,14),
		conv_std_logic_vector(-3677,14),
		conv_std_logic_vector(-3683,14),
		conv_std_logic_vector(-3688,14),
		conv_std_logic_vector(-3694,14),
		conv_std_logic_vector(-3700,14),
		conv_std_logic_vector(-3705,14),
		conv_std_logic_vector(-3711,14),
		conv_std_logic_vector(-3716,14),
		conv_std_logic_vector(-3722,14),
		conv_std_logic_vector(-3728,14),
		conv_std_logic_vector(-3733,14),
		conv_std_logic_vector(-3739,14),
		conv_std_logic_vector(-3744,14),
		conv_std_logic_vector(-3750,14),
		conv_std_logic_vector(-3755,14),
		conv_std_logic_vector(-3761,14),
		conv_std_logic_vector(-3767,14),
		conv_std_logic_vector(-3772,14),
		conv_std_logic_vector(-3778,14),
		conv_std_logic_vector(-3783,14),
		conv_std_logic_vector(-3789,14),
		conv_std_logic_vector(-3795,14),
		conv_std_logic_vector(-3800,14),
		conv_std_logic_vector(-3806,14),
		conv_std_logic_vector(-3811,14),
		conv_std_logic_vector(-3817,14),
		conv_std_logic_vector(-3822,14),
		conv_std_logic_vector(-3828,14),
		conv_std_logic_vector(-3833,14),
		conv_std_logic_vector(-3839,14),
		conv_std_logic_vector(-3845,14),
		conv_std_logic_vector(-3850,14),
		conv_std_logic_vector(-3856,14),
		conv_std_logic_vector(-3861,14),
		conv_std_logic_vector(-3867,14),
		conv_std_logic_vector(-3872,14),
		conv_std_logic_vector(-3878,14),
		conv_std_logic_vector(-3883,14),
		conv_std_logic_vector(-3889,14),
		conv_std_logic_vector(-3894,14),
		conv_std_logic_vector(-3900,14),
		conv_std_logic_vector(-3905,14),
		conv_std_logic_vector(-3911,14),
		conv_std_logic_vector(-3916,14),
		conv_std_logic_vector(-3922,14),
		conv_std_logic_vector(-3928,14),
		conv_std_logic_vector(-3933,14),
		conv_std_logic_vector(-3939,14),
		conv_std_logic_vector(-3944,14),
		conv_std_logic_vector(-3950,14),
		conv_std_logic_vector(-3955,14),
		conv_std_logic_vector(-3961,14),
		conv_std_logic_vector(-3966,14),
		conv_std_logic_vector(-3972,14),
		conv_std_logic_vector(-3977,14),
		conv_std_logic_vector(-3983,14),
		conv_std_logic_vector(-3988,14),
		conv_std_logic_vector(-3994,14),
		conv_std_logic_vector(-3999,14),
		conv_std_logic_vector(-4004,14),
		conv_std_logic_vector(-4010,14),
		conv_std_logic_vector(-4015,14),
		conv_std_logic_vector(-4021,14),
		conv_std_logic_vector(-4026,14),
		conv_std_logic_vector(-4032,14),
		conv_std_logic_vector(-4037,14),
		conv_std_logic_vector(-4043,14),
		conv_std_logic_vector(-4048,14),
		conv_std_logic_vector(-4054,14),
		conv_std_logic_vector(-4059,14),
		conv_std_logic_vector(-4065,14),
		conv_std_logic_vector(-4070,14),
		conv_std_logic_vector(-4076,14),
		conv_std_logic_vector(-4081,14),
		conv_std_logic_vector(-4086,14),
		conv_std_logic_vector(-4092,14),
		conv_std_logic_vector(-4097,14),
		conv_std_logic_vector(-4103,14),
		conv_std_logic_vector(-4108,14),
		conv_std_logic_vector(-4114,14),
		conv_std_logic_vector(-4119,14),
		conv_std_logic_vector(-4124,14),
		conv_std_logic_vector(-4130,14),
		conv_std_logic_vector(-4135,14),
		conv_std_logic_vector(-4141,14),
		conv_std_logic_vector(-4146,14),
		conv_std_logic_vector(-4152,14),
		conv_std_logic_vector(-4157,14),
		conv_std_logic_vector(-4162,14),
		conv_std_logic_vector(-4168,14),
		conv_std_logic_vector(-4173,14),
		conv_std_logic_vector(-4179,14),
		conv_std_logic_vector(-4184,14),
		conv_std_logic_vector(-4189,14),
		conv_std_logic_vector(-4195,14),
		conv_std_logic_vector(-4200,14),
		conv_std_logic_vector(-4206,14),
		conv_std_logic_vector(-4211,14),
		conv_std_logic_vector(-4216,14),
		conv_std_logic_vector(-4222,14),
		conv_std_logic_vector(-4227,14),
		conv_std_logic_vector(-4233,14),
		conv_std_logic_vector(-4238,14),
		conv_std_logic_vector(-4243,14),
		conv_std_logic_vector(-4249,14),
		conv_std_logic_vector(-4254,14),
		conv_std_logic_vector(-4259,14),
		conv_std_logic_vector(-4265,14),
		conv_std_logic_vector(-4270,14),
		conv_std_logic_vector(-4276,14),
		conv_std_logic_vector(-4281,14),
		conv_std_logic_vector(-4286,14),
		conv_std_logic_vector(-4292,14),
		conv_std_logic_vector(-4297,14),
		conv_std_logic_vector(-4302,14),
		conv_std_logic_vector(-4308,14),
		conv_std_logic_vector(-4313,14),
		conv_std_logic_vector(-4318,14),
		conv_std_logic_vector(-4324,14),
		conv_std_logic_vector(-4329,14),
		conv_std_logic_vector(-4334,14),
		conv_std_logic_vector(-4340,14),
		conv_std_logic_vector(-4345,14),
		conv_std_logic_vector(-4350,14),
		conv_std_logic_vector(-4356,14),
		conv_std_logic_vector(-4361,14),
		conv_std_logic_vector(-4366,14),
		conv_std_logic_vector(-4372,14),
		conv_std_logic_vector(-4377,14),
		conv_std_logic_vector(-4382,14),
		conv_std_logic_vector(-4388,14),
		conv_std_logic_vector(-4393,14),
		conv_std_logic_vector(-4398,14),
		conv_std_logic_vector(-4403,14),
		conv_std_logic_vector(-4409,14),
		conv_std_logic_vector(-4414,14),
		conv_std_logic_vector(-4419,14),
		conv_std_logic_vector(-4425,14),
		conv_std_logic_vector(-4430,14),
		conv_std_logic_vector(-4435,14),
		conv_std_logic_vector(-4440,14),
		conv_std_logic_vector(-4446,14),
		conv_std_logic_vector(-4451,14),
		conv_std_logic_vector(-4456,14),
		conv_std_logic_vector(-4462,14),
		conv_std_logic_vector(-4467,14),
		conv_std_logic_vector(-4472,14),
		conv_std_logic_vector(-4477,14),
		conv_std_logic_vector(-4483,14),
		conv_std_logic_vector(-4488,14),
		conv_std_logic_vector(-4493,14),
		conv_std_logic_vector(-4498,14),
		conv_std_logic_vector(-4504,14),
		conv_std_logic_vector(-4509,14),
		conv_std_logic_vector(-4514,14),
		conv_std_logic_vector(-4519,14),
		conv_std_logic_vector(-4525,14),
		conv_std_logic_vector(-4530,14),
		conv_std_logic_vector(-4535,14),
		conv_std_logic_vector(-4540,14),
		conv_std_logic_vector(-4546,14),
		conv_std_logic_vector(-4551,14),
		conv_std_logic_vector(-4556,14),
		conv_std_logic_vector(-4561,14),
		conv_std_logic_vector(-4566,14),
		conv_std_logic_vector(-4572,14),
		conv_std_logic_vector(-4577,14),
		conv_std_logic_vector(-4582,14),
		conv_std_logic_vector(-4587,14),
		conv_std_logic_vector(-4592,14),
		conv_std_logic_vector(-4598,14),
		conv_std_logic_vector(-4603,14),
		conv_std_logic_vector(-4608,14),
		conv_std_logic_vector(-4613,14),
		conv_std_logic_vector(-4618,14),
		conv_std_logic_vector(-4624,14),
		conv_std_logic_vector(-4629,14),
		conv_std_logic_vector(-4634,14),
		conv_std_logic_vector(-4639,14),
		conv_std_logic_vector(-4644,14),
		conv_std_logic_vector(-4650,14),
		conv_std_logic_vector(-4655,14),
		conv_std_logic_vector(-4660,14),
		conv_std_logic_vector(-4665,14),
		conv_std_logic_vector(-4670,14),
		conv_std_logic_vector(-4675,14),
		conv_std_logic_vector(-4680,14),
		conv_std_logic_vector(-4686,14),
		conv_std_logic_vector(-4691,14),
		conv_std_logic_vector(-4696,14),
		conv_std_logic_vector(-4701,14),
		conv_std_logic_vector(-4706,14),
		conv_std_logic_vector(-4711,14),
		conv_std_logic_vector(-4717,14),
		conv_std_logic_vector(-4722,14),
		conv_std_logic_vector(-4727,14),
		conv_std_logic_vector(-4732,14),
		conv_std_logic_vector(-4737,14),
		conv_std_logic_vector(-4742,14),
		conv_std_logic_vector(-4747,14),
		conv_std_logic_vector(-4752,14),
		conv_std_logic_vector(-4758,14),
		conv_std_logic_vector(-4763,14),
		conv_std_logic_vector(-4768,14),
		conv_std_logic_vector(-4773,14),
		conv_std_logic_vector(-4778,14),
		conv_std_logic_vector(-4783,14),
		conv_std_logic_vector(-4788,14),
		conv_std_logic_vector(-4793,14),
		conv_std_logic_vector(-4798,14),
		conv_std_logic_vector(-4803,14),
		conv_std_logic_vector(-4809,14),
		conv_std_logic_vector(-4814,14),
		conv_std_logic_vector(-4819,14),
		conv_std_logic_vector(-4824,14),
		conv_std_logic_vector(-4829,14),
		conv_std_logic_vector(-4834,14),
		conv_std_logic_vector(-4839,14),
		conv_std_logic_vector(-4844,14),
		conv_std_logic_vector(-4849,14),
		conv_std_logic_vector(-4854,14),
		conv_std_logic_vector(-4859,14),
		conv_std_logic_vector(-4864,14),
		conv_std_logic_vector(-4869,14),
		conv_std_logic_vector(-4874,14),
		conv_std_logic_vector(-4879,14),
		conv_std_logic_vector(-4885,14),
		conv_std_logic_vector(-4890,14),
		conv_std_logic_vector(-4895,14),
		conv_std_logic_vector(-4900,14),
		conv_std_logic_vector(-4905,14),
		conv_std_logic_vector(-4910,14),
		conv_std_logic_vector(-4915,14),
		conv_std_logic_vector(-4920,14),
		conv_std_logic_vector(-4925,14),
		conv_std_logic_vector(-4930,14),
		conv_std_logic_vector(-4935,14),
		conv_std_logic_vector(-4940,14),
		conv_std_logic_vector(-4945,14),
		conv_std_logic_vector(-4950,14),
		conv_std_logic_vector(-4955,14),
		conv_std_logic_vector(-4960,14),
		conv_std_logic_vector(-4965,14),
		conv_std_logic_vector(-4970,14),
		conv_std_logic_vector(-4975,14),
		conv_std_logic_vector(-4980,14),
		conv_std_logic_vector(-4985,14),
		conv_std_logic_vector(-4990,14),
		conv_std_logic_vector(-4995,14),
		conv_std_logic_vector(-5000,14),
		conv_std_logic_vector(-5005,14),
		conv_std_logic_vector(-5010,14),
		conv_std_logic_vector(-5015,14),
		conv_std_logic_vector(-5020,14),
		conv_std_logic_vector(-5025,14),
		conv_std_logic_vector(-5030,14),
		conv_std_logic_vector(-5035,14),
		conv_std_logic_vector(-5039,14),
		conv_std_logic_vector(-5044,14),
		conv_std_logic_vector(-5049,14),
		conv_std_logic_vector(-5054,14),
		conv_std_logic_vector(-5059,14),
		conv_std_logic_vector(-5064,14),
		conv_std_logic_vector(-5069,14),
		conv_std_logic_vector(-5074,14),
		conv_std_logic_vector(-5079,14),
		conv_std_logic_vector(-5084,14),
		conv_std_logic_vector(-5089,14),
		conv_std_logic_vector(-5094,14),
		conv_std_logic_vector(-5099,14),
		conv_std_logic_vector(-5104,14),
		conv_std_logic_vector(-5109,14),
		conv_std_logic_vector(-5113,14),
		conv_std_logic_vector(-5118,14),
		conv_std_logic_vector(-5123,14),
		conv_std_logic_vector(-5128,14),
		conv_std_logic_vector(-5133,14),
		conv_std_logic_vector(-5138,14),
		conv_std_logic_vector(-5143,14),
		conv_std_logic_vector(-5148,14),
		conv_std_logic_vector(-5153,14),
		conv_std_logic_vector(-5157,14),
		conv_std_logic_vector(-5162,14),
		conv_std_logic_vector(-5167,14),
		conv_std_logic_vector(-5172,14),
		conv_std_logic_vector(-5177,14),
		conv_std_logic_vector(-5182,14),
		conv_std_logic_vector(-5187,14),
		conv_std_logic_vector(-5192,14),
		conv_std_logic_vector(-5196,14),
		conv_std_logic_vector(-5201,14),
		conv_std_logic_vector(-5206,14),
		conv_std_logic_vector(-5211,14),
		conv_std_logic_vector(-5216,14),
		conv_std_logic_vector(-5221,14),
		conv_std_logic_vector(-5226,14),
		conv_std_logic_vector(-5230,14),
		conv_std_logic_vector(-5235,14),
		conv_std_logic_vector(-5240,14),
		conv_std_logic_vector(-5245,14),
		conv_std_logic_vector(-5250,14),
		conv_std_logic_vector(-5255,14),
		conv_std_logic_vector(-5259,14),
		conv_std_logic_vector(-5264,14),
		conv_std_logic_vector(-5269,14),
		conv_std_logic_vector(-5274,14),
		conv_std_logic_vector(-5279,14),
		conv_std_logic_vector(-5283,14),
		conv_std_logic_vector(-5288,14),
		conv_std_logic_vector(-5293,14),
		conv_std_logic_vector(-5298,14),
		conv_std_logic_vector(-5303,14),
		conv_std_logic_vector(-5307,14),
		conv_std_logic_vector(-5312,14),
		conv_std_logic_vector(-5317,14),
		conv_std_logic_vector(-5322,14),
		conv_std_logic_vector(-5326,14),
		conv_std_logic_vector(-5331,14),
		conv_std_logic_vector(-5336,14),
		conv_std_logic_vector(-5341,14),
		conv_std_logic_vector(-5346,14),
		conv_std_logic_vector(-5350,14),
		conv_std_logic_vector(-5355,14),
		conv_std_logic_vector(-5360,14),
		conv_std_logic_vector(-5365,14),
		conv_std_logic_vector(-5369,14),
		conv_std_logic_vector(-5374,14),
		conv_std_logic_vector(-5379,14),
		conv_std_logic_vector(-5384,14),
		conv_std_logic_vector(-5388,14),
		conv_std_logic_vector(-5393,14),
		conv_std_logic_vector(-5398,14),
		conv_std_logic_vector(-5402,14),
		conv_std_logic_vector(-5407,14),
		conv_std_logic_vector(-5412,14),
		conv_std_logic_vector(-5417,14),
		conv_std_logic_vector(-5421,14),
		conv_std_logic_vector(-5426,14),
		conv_std_logic_vector(-5431,14),
		conv_std_logic_vector(-5435,14),
		conv_std_logic_vector(-5440,14),
		conv_std_logic_vector(-5445,14),
		conv_std_logic_vector(-5450,14),
		conv_std_logic_vector(-5454,14),
		conv_std_logic_vector(-5459,14),
		conv_std_logic_vector(-5464,14),
		conv_std_logic_vector(-5468,14),
		conv_std_logic_vector(-5473,14),
		conv_std_logic_vector(-5478,14),
		conv_std_logic_vector(-5482,14),
		conv_std_logic_vector(-5487,14),
		conv_std_logic_vector(-5492,14),
		conv_std_logic_vector(-5496,14),
		conv_std_logic_vector(-5501,14),
		conv_std_logic_vector(-5506,14),
		conv_std_logic_vector(-5510,14),
		conv_std_logic_vector(-5515,14),
		conv_std_logic_vector(-5520,14),
		conv_std_logic_vector(-5524,14),
		conv_std_logic_vector(-5529,14),
		conv_std_logic_vector(-5533,14),
		conv_std_logic_vector(-5538,14),
		conv_std_logic_vector(-5543,14),
		conv_std_logic_vector(-5547,14),
		conv_std_logic_vector(-5552,14),
		conv_std_logic_vector(-5557,14),
		conv_std_logic_vector(-5561,14),
		conv_std_logic_vector(-5566,14),
		conv_std_logic_vector(-5570,14),
		conv_std_logic_vector(-5575,14),
		conv_std_logic_vector(-5580,14),
		conv_std_logic_vector(-5584,14),
		conv_std_logic_vector(-5589,14),
		conv_std_logic_vector(-5593,14),
		conv_std_logic_vector(-5598,14),
		conv_std_logic_vector(-5603,14),
		conv_std_logic_vector(-5607,14),
		conv_std_logic_vector(-5612,14),
		conv_std_logic_vector(-5616,14),
		conv_std_logic_vector(-5621,14),
		conv_std_logic_vector(-5625,14),
		conv_std_logic_vector(-5630,14),
		conv_std_logic_vector(-5635,14),
		conv_std_logic_vector(-5639,14),
		conv_std_logic_vector(-5644,14),
		conv_std_logic_vector(-5648,14),
		conv_std_logic_vector(-5653,14),
		conv_std_logic_vector(-5657,14),
		conv_std_logic_vector(-5662,14),
		conv_std_logic_vector(-5666,14),
		conv_std_logic_vector(-5671,14),
		conv_std_logic_vector(-5675,14),
		conv_std_logic_vector(-5680,14),
		conv_std_logic_vector(-5685,14),
		conv_std_logic_vector(-5689,14),
		conv_std_logic_vector(-5694,14),
		conv_std_logic_vector(-5698,14),
		conv_std_logic_vector(-5703,14),
		conv_std_logic_vector(-5707,14),
		conv_std_logic_vector(-5712,14),
		conv_std_logic_vector(-5716,14),
		conv_std_logic_vector(-5721,14),
		conv_std_logic_vector(-5725,14),
		conv_std_logic_vector(-5730,14),
		conv_std_logic_vector(-5734,14),
		conv_std_logic_vector(-5739,14),
		conv_std_logic_vector(-5743,14),
		conv_std_logic_vector(-5748,14),
		conv_std_logic_vector(-5752,14),
		conv_std_logic_vector(-5756,14),
		conv_std_logic_vector(-5761,14),
		conv_std_logic_vector(-5765,14),
		conv_std_logic_vector(-5770,14),
		conv_std_logic_vector(-5774,14),
		conv_std_logic_vector(-5779,14),
		conv_std_logic_vector(-5783,14),
		conv_std_logic_vector(-5788,14),
		conv_std_logic_vector(-5792,14),
		conv_std_logic_vector(-5797,14),
		conv_std_logic_vector(-5801,14),
		conv_std_logic_vector(-5805,14),
		conv_std_logic_vector(-5810,14),
		conv_std_logic_vector(-5814,14),
		conv_std_logic_vector(-5819,14),
		conv_std_logic_vector(-5823,14),
		conv_std_logic_vector(-5828,14),
		conv_std_logic_vector(-5832,14),
		conv_std_logic_vector(-5836,14),
		conv_std_logic_vector(-5841,14),
		conv_std_logic_vector(-5845,14),
		conv_std_logic_vector(-5850,14),
		conv_std_logic_vector(-5854,14),
		conv_std_logic_vector(-5858,14),
		conv_std_logic_vector(-5863,14),
		conv_std_logic_vector(-5867,14),
		conv_std_logic_vector(-5872,14),
		conv_std_logic_vector(-5876,14),
		conv_std_logic_vector(-5880,14),
		conv_std_logic_vector(-5885,14),
		conv_std_logic_vector(-5889,14),
		conv_std_logic_vector(-5893,14),
		conv_std_logic_vector(-5898,14),
		conv_std_logic_vector(-5902,14),
		conv_std_logic_vector(-5906,14),
		conv_std_logic_vector(-5911,14),
		conv_std_logic_vector(-5915,14),
		conv_std_logic_vector(-5920,14),
		conv_std_logic_vector(-5924,14),
		conv_std_logic_vector(-5928,14),
		conv_std_logic_vector(-5933,14),
		conv_std_logic_vector(-5937,14),
		conv_std_logic_vector(-5941,14),
		conv_std_logic_vector(-5946,14),
		conv_std_logic_vector(-5950,14),
		conv_std_logic_vector(-5954,14),
		conv_std_logic_vector(-5958,14),
		conv_std_logic_vector(-5963,14),
		conv_std_logic_vector(-5967,14),
		conv_std_logic_vector(-5971,14),
		conv_std_logic_vector(-5976,14),
		conv_std_logic_vector(-5980,14),
		conv_std_logic_vector(-5984,14),
		conv_std_logic_vector(-5989,14),
		conv_std_logic_vector(-5993,14),
		conv_std_logic_vector(-5997,14),
		conv_std_logic_vector(-6001,14),
		conv_std_logic_vector(-6006,14),
		conv_std_logic_vector(-6010,14),
		conv_std_logic_vector(-6014,14),
		conv_std_logic_vector(-6018,14),
		conv_std_logic_vector(-6023,14),
		conv_std_logic_vector(-6027,14),
		conv_std_logic_vector(-6031,14),
		conv_std_logic_vector(-6036,14),
		conv_std_logic_vector(-6040,14),
		conv_std_logic_vector(-6044,14),
		conv_std_logic_vector(-6048,14),
		conv_std_logic_vector(-6052,14),
		conv_std_logic_vector(-6057,14),
		conv_std_logic_vector(-6061,14),
		conv_std_logic_vector(-6065,14),
		conv_std_logic_vector(-6069,14),
		conv_std_logic_vector(-6074,14),
		conv_std_logic_vector(-6078,14),
		conv_std_logic_vector(-6082,14),
		conv_std_logic_vector(-6086,14),
		conv_std_logic_vector(-6090,14),
		conv_std_logic_vector(-6095,14),
		conv_std_logic_vector(-6099,14),
		conv_std_logic_vector(-6103,14),
		conv_std_logic_vector(-6107,14),
		conv_std_logic_vector(-6111,14),
		conv_std_logic_vector(-6116,14),
		conv_std_logic_vector(-6120,14),
		conv_std_logic_vector(-6124,14),
		conv_std_logic_vector(-6128,14),
		conv_std_logic_vector(-6132,14),
		conv_std_logic_vector(-6136,14),
		conv_std_logic_vector(-6141,14),
		conv_std_logic_vector(-6145,14),
		conv_std_logic_vector(-6149,14),
		conv_std_logic_vector(-6153,14),
		conv_std_logic_vector(-6157,14),
		conv_std_logic_vector(-6161,14),
		conv_std_logic_vector(-6165,14),
		conv_std_logic_vector(-6170,14),
		conv_std_logic_vector(-6174,14),
		conv_std_logic_vector(-6178,14),
		conv_std_logic_vector(-6182,14),
		conv_std_logic_vector(-6186,14),
		conv_std_logic_vector(-6190,14),
		conv_std_logic_vector(-6194,14),
		conv_std_logic_vector(-6198,14),
		conv_std_logic_vector(-6203,14),
		conv_std_logic_vector(-6207,14),
		conv_std_logic_vector(-6211,14),
		conv_std_logic_vector(-6215,14),
		conv_std_logic_vector(-6219,14),
		conv_std_logic_vector(-6223,14),
		conv_std_logic_vector(-6227,14),
		conv_std_logic_vector(-6231,14),
		conv_std_logic_vector(-6235,14),
		conv_std_logic_vector(-6239,14),
		conv_std_logic_vector(-6243,14),
		conv_std_logic_vector(-6247,14),
		conv_std_logic_vector(-6252,14),
		conv_std_logic_vector(-6256,14),
		conv_std_logic_vector(-6260,14),
		conv_std_logic_vector(-6264,14),
		conv_std_logic_vector(-6268,14),
		conv_std_logic_vector(-6272,14),
		conv_std_logic_vector(-6276,14),
		conv_std_logic_vector(-6280,14),
		conv_std_logic_vector(-6284,14),
		conv_std_logic_vector(-6288,14),
		conv_std_logic_vector(-6292,14),
		conv_std_logic_vector(-6296,14),
		conv_std_logic_vector(-6300,14),
		conv_std_logic_vector(-6304,14),
		conv_std_logic_vector(-6308,14),
		conv_std_logic_vector(-6312,14),
		conv_std_logic_vector(-6316,14),
		conv_std_logic_vector(-6320,14),
		conv_std_logic_vector(-6324,14),
		conv_std_logic_vector(-6328,14),
		conv_std_logic_vector(-6332,14),
		conv_std_logic_vector(-6336,14),
		conv_std_logic_vector(-6340,14),
		conv_std_logic_vector(-6344,14),
		conv_std_logic_vector(-6348,14),
		conv_std_logic_vector(-6352,14),
		conv_std_logic_vector(-6356,14),
		conv_std_logic_vector(-6360,14),
		conv_std_logic_vector(-6364,14),
		conv_std_logic_vector(-6368,14),
		conv_std_logic_vector(-6372,14),
		conv_std_logic_vector(-6376,14),
		conv_std_logic_vector(-6380,14),
		conv_std_logic_vector(-6384,14),
		conv_std_logic_vector(-6387,14),
		conv_std_logic_vector(-6391,14),
		conv_std_logic_vector(-6395,14),
		conv_std_logic_vector(-6399,14),
		conv_std_logic_vector(-6403,14),
		conv_std_logic_vector(-6407,14),
		conv_std_logic_vector(-6411,14),
		conv_std_logic_vector(-6415,14),
		conv_std_logic_vector(-6419,14),
		conv_std_logic_vector(-6423,14),
		conv_std_logic_vector(-6427,14),
		conv_std_logic_vector(-6430,14),
		conv_std_logic_vector(-6434,14),
		conv_std_logic_vector(-6438,14),
		conv_std_logic_vector(-6442,14),
		conv_std_logic_vector(-6446,14),
		conv_std_logic_vector(-6450,14),
		conv_std_logic_vector(-6454,14),
		conv_std_logic_vector(-6458,14),
		conv_std_logic_vector(-6461,14),
		conv_std_logic_vector(-6465,14),
		conv_std_logic_vector(-6469,14),
		conv_std_logic_vector(-6473,14),
		conv_std_logic_vector(-6477,14),
		conv_std_logic_vector(-6481,14),
		conv_std_logic_vector(-6485,14),
		conv_std_logic_vector(-6488,14),
		conv_std_logic_vector(-6492,14),
		conv_std_logic_vector(-6496,14),
		conv_std_logic_vector(-6500,14),
		conv_std_logic_vector(-6504,14),
		conv_std_logic_vector(-6508,14),
		conv_std_logic_vector(-6511,14),
		conv_std_logic_vector(-6515,14),
		conv_std_logic_vector(-6519,14),
		conv_std_logic_vector(-6523,14),
		conv_std_logic_vector(-6527,14),
		conv_std_logic_vector(-6530,14),
		conv_std_logic_vector(-6534,14),
		conv_std_logic_vector(-6538,14),
		conv_std_logic_vector(-6542,14),
		conv_std_logic_vector(-6546,14),
		conv_std_logic_vector(-6549,14),
		conv_std_logic_vector(-6553,14),
		conv_std_logic_vector(-6557,14),
		conv_std_logic_vector(-6561,14),
		conv_std_logic_vector(-6564,14),
		conv_std_logic_vector(-6568,14),
		conv_std_logic_vector(-6572,14),
		conv_std_logic_vector(-6576,14),
		conv_std_logic_vector(-6579,14),
		conv_std_logic_vector(-6583,14),
		conv_std_logic_vector(-6587,14),
		conv_std_logic_vector(-6591,14),
		conv_std_logic_vector(-6594,14),
		conv_std_logic_vector(-6598,14),
		conv_std_logic_vector(-6602,14),
		conv_std_logic_vector(-6605,14),
		conv_std_logic_vector(-6609,14),
		conv_std_logic_vector(-6613,14),
		conv_std_logic_vector(-6617,14),
		conv_std_logic_vector(-6620,14),
		conv_std_logic_vector(-6624,14),
		conv_std_logic_vector(-6628,14),
		conv_std_logic_vector(-6631,14),
		conv_std_logic_vector(-6635,14),
		conv_std_logic_vector(-6639,14),
		conv_std_logic_vector(-6642,14),
		conv_std_logic_vector(-6646,14),
		conv_std_logic_vector(-6650,14),
		conv_std_logic_vector(-6653,14),
		conv_std_logic_vector(-6657,14),
		conv_std_logic_vector(-6661,14),
		conv_std_logic_vector(-6664,14),
		conv_std_logic_vector(-6668,14),
		conv_std_logic_vector(-6672,14),
		conv_std_logic_vector(-6675,14),
		conv_std_logic_vector(-6679,14),
		conv_std_logic_vector(-6683,14),
		conv_std_logic_vector(-6686,14),
		conv_std_logic_vector(-6690,14),
		conv_std_logic_vector(-6694,14),
		conv_std_logic_vector(-6697,14),
		conv_std_logic_vector(-6701,14),
		conv_std_logic_vector(-6704,14),
		conv_std_logic_vector(-6708,14),
		conv_std_logic_vector(-6712,14),
		conv_std_logic_vector(-6715,14),
		conv_std_logic_vector(-6719,14),
		conv_std_logic_vector(-6722,14),
		conv_std_logic_vector(-6726,14),
		conv_std_logic_vector(-6730,14),
		conv_std_logic_vector(-6733,14),
		conv_std_logic_vector(-6737,14),
		conv_std_logic_vector(-6740,14),
		conv_std_logic_vector(-6744,14),
		conv_std_logic_vector(-6747,14),
		conv_std_logic_vector(-6751,14),
		conv_std_logic_vector(-6755,14),
		conv_std_logic_vector(-6758,14),
		conv_std_logic_vector(-6762,14),
		conv_std_logic_vector(-6765,14),
		conv_std_logic_vector(-6769,14),
		conv_std_logic_vector(-6772,14),
		conv_std_logic_vector(-6776,14),
		conv_std_logic_vector(-6779,14),
		conv_std_logic_vector(-6783,14),
		conv_std_logic_vector(-6786,14),
		conv_std_logic_vector(-6790,14),
		conv_std_logic_vector(-6793,14),
		conv_std_logic_vector(-6797,14),
		conv_std_logic_vector(-6800,14),
		conv_std_logic_vector(-6804,14),
		conv_std_logic_vector(-6807,14),
		conv_std_logic_vector(-6811,14),
		conv_std_logic_vector(-6814,14),
		conv_std_logic_vector(-6818,14),
		conv_std_logic_vector(-6821,14),
		conv_std_logic_vector(-6825,14),
		conv_std_logic_vector(-6828,14),
		conv_std_logic_vector(-6832,14),
		conv_std_logic_vector(-6835,14),
		conv_std_logic_vector(-6839,14),
		conv_std_logic_vector(-6842,14),
		conv_std_logic_vector(-6846,14),
		conv_std_logic_vector(-6849,14),
		conv_std_logic_vector(-6852,14),
		conv_std_logic_vector(-6856,14),
		conv_std_logic_vector(-6859,14),
		conv_std_logic_vector(-6863,14),
		conv_std_logic_vector(-6866,14),
		conv_std_logic_vector(-6870,14),
		conv_std_logic_vector(-6873,14),
		conv_std_logic_vector(-6876,14),
		conv_std_logic_vector(-6880,14),
		conv_std_logic_vector(-6883,14),
		conv_std_logic_vector(-6887,14),
		conv_std_logic_vector(-6890,14),
		conv_std_logic_vector(-6894,14),
		conv_std_logic_vector(-6897,14),
		conv_std_logic_vector(-6900,14),
		conv_std_logic_vector(-6904,14),
		conv_std_logic_vector(-6907,14),
		conv_std_logic_vector(-6910,14),
		conv_std_logic_vector(-6914,14),
		conv_std_logic_vector(-6917,14),
		conv_std_logic_vector(-6921,14),
		conv_std_logic_vector(-6924,14),
		conv_std_logic_vector(-6927,14),
		conv_std_logic_vector(-6931,14),
		conv_std_logic_vector(-6934,14),
		conv_std_logic_vector(-6937,14),
		conv_std_logic_vector(-6941,14),
		conv_std_logic_vector(-6944,14),
		conv_std_logic_vector(-6947,14),
		conv_std_logic_vector(-6951,14),
		conv_std_logic_vector(-6954,14),
		conv_std_logic_vector(-6957,14),
		conv_std_logic_vector(-6961,14),
		conv_std_logic_vector(-6964,14),
		conv_std_logic_vector(-6967,14),
		conv_std_logic_vector(-6971,14),
		conv_std_logic_vector(-6974,14),
		conv_std_logic_vector(-6977,14),
		conv_std_logic_vector(-6980,14),
		conv_std_logic_vector(-6984,14),
		conv_std_logic_vector(-6987,14),
		conv_std_logic_vector(-6990,14),
		conv_std_logic_vector(-6994,14),
		conv_std_logic_vector(-6997,14),
		conv_std_logic_vector(-7000,14),
		conv_std_logic_vector(-7003,14),
		conv_std_logic_vector(-7007,14),
		conv_std_logic_vector(-7010,14),
		conv_std_logic_vector(-7013,14),
		conv_std_logic_vector(-7016,14),
		conv_std_logic_vector(-7020,14),
		conv_std_logic_vector(-7023,14),
		conv_std_logic_vector(-7026,14),
		conv_std_logic_vector(-7029,14),
		conv_std_logic_vector(-7032,14),
		conv_std_logic_vector(-7036,14),
		conv_std_logic_vector(-7039,14),
		conv_std_logic_vector(-7042,14),
		conv_std_logic_vector(-7045,14),
		conv_std_logic_vector(-7049,14),
		conv_std_logic_vector(-7052,14),
		conv_std_logic_vector(-7055,14),
		conv_std_logic_vector(-7058,14),
		conv_std_logic_vector(-7061,14),
		conv_std_logic_vector(-7064,14),
		conv_std_logic_vector(-7068,14),
		conv_std_logic_vector(-7071,14),
		conv_std_logic_vector(-7074,14),
		conv_std_logic_vector(-7077,14),
		conv_std_logic_vector(-7080,14),
		conv_std_logic_vector(-7083,14),
		conv_std_logic_vector(-7087,14),
		conv_std_logic_vector(-7090,14),
		conv_std_logic_vector(-7093,14),
		conv_std_logic_vector(-7096,14),
		conv_std_logic_vector(-7099,14),
		conv_std_logic_vector(-7102,14),
		conv_std_logic_vector(-7105,14),
		conv_std_logic_vector(-7109,14),
		conv_std_logic_vector(-7112,14),
		conv_std_logic_vector(-7115,14),
		conv_std_logic_vector(-7118,14),
		conv_std_logic_vector(-7121,14),
		conv_std_logic_vector(-7124,14),
		conv_std_logic_vector(-7127,14),
		conv_std_logic_vector(-7130,14),
		conv_std_logic_vector(-7133,14),
		conv_std_logic_vector(-7137,14),
		conv_std_logic_vector(-7140,14),
		conv_std_logic_vector(-7143,14),
		conv_std_logic_vector(-7146,14),
		conv_std_logic_vector(-7149,14),
		conv_std_logic_vector(-7152,14),
		conv_std_logic_vector(-7155,14),
		conv_std_logic_vector(-7158,14),
		conv_std_logic_vector(-7161,14),
		conv_std_logic_vector(-7164,14),
		conv_std_logic_vector(-7167,14),
		conv_std_logic_vector(-7170,14),
		conv_std_logic_vector(-7173,14),
		conv_std_logic_vector(-7176,14),
		conv_std_logic_vector(-7179,14),
		conv_std_logic_vector(-7182,14),
		conv_std_logic_vector(-7185,14),
		conv_std_logic_vector(-7188,14),
		conv_std_logic_vector(-7191,14),
		conv_std_logic_vector(-7194,14),
		conv_std_logic_vector(-7197,14),
		conv_std_logic_vector(-7200,14),
		conv_std_logic_vector(-7203,14),
		conv_std_logic_vector(-7206,14),
		conv_std_logic_vector(-7209,14),
		conv_std_logic_vector(-7212,14),
		conv_std_logic_vector(-7215,14),
		conv_std_logic_vector(-7218,14),
		conv_std_logic_vector(-7221,14),
		conv_std_logic_vector(-7224,14),
		conv_std_logic_vector(-7227,14),
		conv_std_logic_vector(-7230,14),
		conv_std_logic_vector(-7233,14),
		conv_std_logic_vector(-7236,14),
		conv_std_logic_vector(-7239,14),
		conv_std_logic_vector(-7242,14),
		conv_std_logic_vector(-7245,14),
		conv_std_logic_vector(-7248,14),
		conv_std_logic_vector(-7251,14),
		conv_std_logic_vector(-7254,14),
		conv_std_logic_vector(-7257,14),
		conv_std_logic_vector(-7259,14),
		conv_std_logic_vector(-7262,14),
		conv_std_logic_vector(-7265,14),
		conv_std_logic_vector(-7268,14),
		conv_std_logic_vector(-7271,14),
		conv_std_logic_vector(-7274,14),
		conv_std_logic_vector(-7277,14),
		conv_std_logic_vector(-7280,14),
		conv_std_logic_vector(-7283,14),
		conv_std_logic_vector(-7285,14),
		conv_std_logic_vector(-7288,14),
		conv_std_logic_vector(-7291,14),
		conv_std_logic_vector(-7294,14),
		conv_std_logic_vector(-7297,14),
		conv_std_logic_vector(-7300,14),
		conv_std_logic_vector(-7303,14),
		conv_std_logic_vector(-7305,14),
		conv_std_logic_vector(-7308,14),
		conv_std_logic_vector(-7311,14),
		conv_std_logic_vector(-7314,14),
		conv_std_logic_vector(-7317,14),
		conv_std_logic_vector(-7320,14),
		conv_std_logic_vector(-7322,14),
		conv_std_logic_vector(-7325,14),
		conv_std_logic_vector(-7328,14),
		conv_std_logic_vector(-7331,14),
		conv_std_logic_vector(-7334,14),
		conv_std_logic_vector(-7336,14),
		conv_std_logic_vector(-7339,14),
		conv_std_logic_vector(-7342,14),
		conv_std_logic_vector(-7345,14),
		conv_std_logic_vector(-7348,14),
		conv_std_logic_vector(-7350,14),
		conv_std_logic_vector(-7353,14),
		conv_std_logic_vector(-7356,14),
		conv_std_logic_vector(-7359,14),
		conv_std_logic_vector(-7361,14),
		conv_std_logic_vector(-7364,14),
		conv_std_logic_vector(-7367,14),
		conv_std_logic_vector(-7370,14),
		conv_std_logic_vector(-7372,14),
		conv_std_logic_vector(-7375,14),
		conv_std_logic_vector(-7378,14),
		conv_std_logic_vector(-7381,14),
		conv_std_logic_vector(-7383,14),
		conv_std_logic_vector(-7386,14),
		conv_std_logic_vector(-7389,14),
		conv_std_logic_vector(-7391,14),
		conv_std_logic_vector(-7394,14),
		conv_std_logic_vector(-7397,14),
		conv_std_logic_vector(-7400,14),
		conv_std_logic_vector(-7402,14),
		conv_std_logic_vector(-7405,14),
		conv_std_logic_vector(-7408,14),
		conv_std_logic_vector(-7410,14),
		conv_std_logic_vector(-7413,14),
		conv_std_logic_vector(-7416,14),
		conv_std_logic_vector(-7418,14),
		conv_std_logic_vector(-7421,14),
		conv_std_logic_vector(-7424,14),
		conv_std_logic_vector(-7426,14),
		conv_std_logic_vector(-7429,14),
		conv_std_logic_vector(-7432,14),
		conv_std_logic_vector(-7434,14),
		conv_std_logic_vector(-7437,14),
		conv_std_logic_vector(-7440,14),
		conv_std_logic_vector(-7442,14),
		conv_std_logic_vector(-7445,14),
		conv_std_logic_vector(-7447,14),
		conv_std_logic_vector(-7450,14),
		conv_std_logic_vector(-7453,14),
		conv_std_logic_vector(-7455,14),
		conv_std_logic_vector(-7458,14),
		conv_std_logic_vector(-7460,14),
		conv_std_logic_vector(-7463,14),
		conv_std_logic_vector(-7466,14),
		conv_std_logic_vector(-7468,14),
		conv_std_logic_vector(-7471,14),
		conv_std_logic_vector(-7473,14),
		conv_std_logic_vector(-7476,14),
		conv_std_logic_vector(-7478,14),
		conv_std_logic_vector(-7481,14),
		conv_std_logic_vector(-7484,14),
		conv_std_logic_vector(-7486,14),
		conv_std_logic_vector(-7489,14),
		conv_std_logic_vector(-7491,14),
		conv_std_logic_vector(-7494,14),
		conv_std_logic_vector(-7496,14),
		conv_std_logic_vector(-7499,14),
		conv_std_logic_vector(-7501,14),
		conv_std_logic_vector(-7504,14),
		conv_std_logic_vector(-7506,14),
		conv_std_logic_vector(-7509,14),
		conv_std_logic_vector(-7511,14),
		conv_std_logic_vector(-7514,14),
		conv_std_logic_vector(-7516,14),
		conv_std_logic_vector(-7519,14),
		conv_std_logic_vector(-7521,14),
		conv_std_logic_vector(-7524,14),
		conv_std_logic_vector(-7526,14),
		conv_std_logic_vector(-7529,14),
		conv_std_logic_vector(-7531,14),
		conv_std_logic_vector(-7534,14),
		conv_std_logic_vector(-7536,14),
		conv_std_logic_vector(-7539,14),
		conv_std_logic_vector(-7541,14),
		conv_std_logic_vector(-7544,14),
		conv_std_logic_vector(-7546,14),
		conv_std_logic_vector(-7549,14),
		conv_std_logic_vector(-7551,14),
		conv_std_logic_vector(-7553,14),
		conv_std_logic_vector(-7556,14),
		conv_std_logic_vector(-7558,14),
		conv_std_logic_vector(-7561,14),
		conv_std_logic_vector(-7563,14),
		conv_std_logic_vector(-7566,14),
		conv_std_logic_vector(-7568,14),
		conv_std_logic_vector(-7570,14),
		conv_std_logic_vector(-7573,14),
		conv_std_logic_vector(-7575,14),
		conv_std_logic_vector(-7578,14),
		conv_std_logic_vector(-7580,14),
		conv_std_logic_vector(-7582,14),
		conv_std_logic_vector(-7585,14),
		conv_std_logic_vector(-7587,14),
		conv_std_logic_vector(-7589,14),
		conv_std_logic_vector(-7592,14),
		conv_std_logic_vector(-7594,14),
		conv_std_logic_vector(-7596,14),
		conv_std_logic_vector(-7599,14),
		conv_std_logic_vector(-7601,14),
		conv_std_logic_vector(-7603,14),
		conv_std_logic_vector(-7606,14),
		conv_std_logic_vector(-7608,14),
		conv_std_logic_vector(-7610,14),
		conv_std_logic_vector(-7613,14),
		conv_std_logic_vector(-7615,14),
		conv_std_logic_vector(-7617,14),
		conv_std_logic_vector(-7620,14),
		conv_std_logic_vector(-7622,14),
		conv_std_logic_vector(-7624,14),
		conv_std_logic_vector(-7627,14),
		conv_std_logic_vector(-7629,14),
		conv_std_logic_vector(-7631,14),
		conv_std_logic_vector(-7633,14),
		conv_std_logic_vector(-7636,14),
		conv_std_logic_vector(-7638,14),
		conv_std_logic_vector(-7640,14),
		conv_std_logic_vector(-7643,14),
		conv_std_logic_vector(-7645,14),
		conv_std_logic_vector(-7647,14),
		conv_std_logic_vector(-7649,14),
		conv_std_logic_vector(-7652,14),
		conv_std_logic_vector(-7654,14),
		conv_std_logic_vector(-7656,14),
		conv_std_logic_vector(-7658,14),
		conv_std_logic_vector(-7661,14),
		conv_std_logic_vector(-7663,14),
		conv_std_logic_vector(-7665,14),
		conv_std_logic_vector(-7667,14),
		conv_std_logic_vector(-7669,14),
		conv_std_logic_vector(-7672,14),
		conv_std_logic_vector(-7674,14),
		conv_std_logic_vector(-7676,14),
		conv_std_logic_vector(-7678,14),
		conv_std_logic_vector(-7680,14),
		conv_std_logic_vector(-7683,14),
		conv_std_logic_vector(-7685,14),
		conv_std_logic_vector(-7687,14),
		conv_std_logic_vector(-7689,14),
		conv_std_logic_vector(-7691,14),
		conv_std_logic_vector(-7693,14),
		conv_std_logic_vector(-7696,14),
		conv_std_logic_vector(-7698,14),
		conv_std_logic_vector(-7700,14),
		conv_std_logic_vector(-7702,14),
		conv_std_logic_vector(-7704,14),
		conv_std_logic_vector(-7706,14),
		conv_std_logic_vector(-7708,14),
		conv_std_logic_vector(-7711,14),
		conv_std_logic_vector(-7713,14),
		conv_std_logic_vector(-7715,14),
		conv_std_logic_vector(-7717,14),
		conv_std_logic_vector(-7719,14),
		conv_std_logic_vector(-7721,14),
		conv_std_logic_vector(-7723,14),
		conv_std_logic_vector(-7725,14),
		conv_std_logic_vector(-7727,14),
		conv_std_logic_vector(-7729,14),
		conv_std_logic_vector(-7731,14),
		conv_std_logic_vector(-7734,14),
		conv_std_logic_vector(-7736,14),
		conv_std_logic_vector(-7738,14),
		conv_std_logic_vector(-7740,14),
		conv_std_logic_vector(-7742,14),
		conv_std_logic_vector(-7744,14),
		conv_std_logic_vector(-7746,14),
		conv_std_logic_vector(-7748,14),
		conv_std_logic_vector(-7750,14),
		conv_std_logic_vector(-7752,14),
		conv_std_logic_vector(-7754,14),
		conv_std_logic_vector(-7756,14),
		conv_std_logic_vector(-7758,14),
		conv_std_logic_vector(-7760,14),
		conv_std_logic_vector(-7762,14),
		conv_std_logic_vector(-7764,14),
		conv_std_logic_vector(-7766,14),
		conv_std_logic_vector(-7768,14),
		conv_std_logic_vector(-7770,14),
		conv_std_logic_vector(-7772,14),
		conv_std_logic_vector(-7774,14),
		conv_std_logic_vector(-7776,14),
		conv_std_logic_vector(-7778,14),
		conv_std_logic_vector(-7780,14),
		conv_std_logic_vector(-7782,14),
		conv_std_logic_vector(-7784,14),
		conv_std_logic_vector(-7786,14),
		conv_std_logic_vector(-7788,14),
		conv_std_logic_vector(-7790,14),
		conv_std_logic_vector(-7792,14),
		conv_std_logic_vector(-7794,14),
		conv_std_logic_vector(-7796,14),
		conv_std_logic_vector(-7798,14),
		conv_std_logic_vector(-7799,14),
		conv_std_logic_vector(-7801,14),
		conv_std_logic_vector(-7803,14),
		conv_std_logic_vector(-7805,14),
		conv_std_logic_vector(-7807,14),
		conv_std_logic_vector(-7809,14),
		conv_std_logic_vector(-7811,14),
		conv_std_logic_vector(-7813,14),
		conv_std_logic_vector(-7815,14),
		conv_std_logic_vector(-7817,14),
		conv_std_logic_vector(-7818,14),
		conv_std_logic_vector(-7820,14),
		conv_std_logic_vector(-7822,14),
		conv_std_logic_vector(-7824,14),
		conv_std_logic_vector(-7826,14),
		conv_std_logic_vector(-7828,14),
		conv_std_logic_vector(-7830,14),
		conv_std_logic_vector(-7831,14),
		conv_std_logic_vector(-7833,14),
		conv_std_logic_vector(-7835,14),
		conv_std_logic_vector(-7837,14),
		conv_std_logic_vector(-7839,14),
		conv_std_logic_vector(-7841,14),
		conv_std_logic_vector(-7842,14),
		conv_std_logic_vector(-7844,14),
		conv_std_logic_vector(-7846,14),
		conv_std_logic_vector(-7848,14),
		conv_std_logic_vector(-7850,14),
		conv_std_logic_vector(-7851,14),
		conv_std_logic_vector(-7853,14),
		conv_std_logic_vector(-7855,14),
		conv_std_logic_vector(-7857,14),
		conv_std_logic_vector(-7859,14),
		conv_std_logic_vector(-7860,14),
		conv_std_logic_vector(-7862,14),
		conv_std_logic_vector(-7864,14),
		conv_std_logic_vector(-7866,14),
		conv_std_logic_vector(-7867,14),
		conv_std_logic_vector(-7869,14),
		conv_std_logic_vector(-7871,14),
		conv_std_logic_vector(-7873,14),
		conv_std_logic_vector(-7874,14),
		conv_std_logic_vector(-7876,14),
		conv_std_logic_vector(-7878,14),
		conv_std_logic_vector(-7879,14),
		conv_std_logic_vector(-7881,14),
		conv_std_logic_vector(-7883,14),
		conv_std_logic_vector(-7885,14),
		conv_std_logic_vector(-7886,14),
		conv_std_logic_vector(-7888,14),
		conv_std_logic_vector(-7890,14),
		conv_std_logic_vector(-7891,14),
		conv_std_logic_vector(-7893,14),
		conv_std_logic_vector(-7895,14),
		conv_std_logic_vector(-7896,14),
		conv_std_logic_vector(-7898,14),
		conv_std_logic_vector(-7900,14),
		conv_std_logic_vector(-7901,14),
		conv_std_logic_vector(-7903,14),
		conv_std_logic_vector(-7905,14),
		conv_std_logic_vector(-7906,14),
		conv_std_logic_vector(-7908,14),
		conv_std_logic_vector(-7910,14),
		conv_std_logic_vector(-7911,14),
		conv_std_logic_vector(-7913,14),
		conv_std_logic_vector(-7915,14),
		conv_std_logic_vector(-7916,14),
		conv_std_logic_vector(-7918,14),
		conv_std_logic_vector(-7919,14),
		conv_std_logic_vector(-7921,14),
		conv_std_logic_vector(-7923,14),
		conv_std_logic_vector(-7924,14),
		conv_std_logic_vector(-7926,14),
		conv_std_logic_vector(-7927,14),
		conv_std_logic_vector(-7929,14),
		conv_std_logic_vector(-7930,14),
		conv_std_logic_vector(-7932,14),
		conv_std_logic_vector(-7934,14),
		conv_std_logic_vector(-7935,14),
		conv_std_logic_vector(-7937,14),
		conv_std_logic_vector(-7938,14),
		conv_std_logic_vector(-7940,14),
		conv_std_logic_vector(-7941,14),
		conv_std_logic_vector(-7943,14),
		conv_std_logic_vector(-7944,14),
		conv_std_logic_vector(-7946,14),
		conv_std_logic_vector(-7948,14),
		conv_std_logic_vector(-7949,14),
		conv_std_logic_vector(-7951,14),
		conv_std_logic_vector(-7952,14),
		conv_std_logic_vector(-7954,14),
		conv_std_logic_vector(-7955,14),
		conv_std_logic_vector(-7957,14),
		conv_std_logic_vector(-7958,14),
		conv_std_logic_vector(-7960,14),
		conv_std_logic_vector(-7961,14),
		conv_std_logic_vector(-7963,14),
		conv_std_logic_vector(-7964,14),
		conv_std_logic_vector(-7965,14),
		conv_std_logic_vector(-7967,14),
		conv_std_logic_vector(-7968,14),
		conv_std_logic_vector(-7970,14),
		conv_std_logic_vector(-7971,14),
		conv_std_logic_vector(-7973,14),
		conv_std_logic_vector(-7974,14),
		conv_std_logic_vector(-7976,14),
		conv_std_logic_vector(-7977,14),
		conv_std_logic_vector(-7978,14),
		conv_std_logic_vector(-7980,14),
		conv_std_logic_vector(-7981,14),
		conv_std_logic_vector(-7983,14),
		conv_std_logic_vector(-7984,14),
		conv_std_logic_vector(-7986,14),
		conv_std_logic_vector(-7987,14),
		conv_std_logic_vector(-7988,14),
		conv_std_logic_vector(-7990,14),
		conv_std_logic_vector(-7991,14),
		conv_std_logic_vector(-7992,14),
		conv_std_logic_vector(-7994,14),
		conv_std_logic_vector(-7995,14),
		conv_std_logic_vector(-7997,14),
		conv_std_logic_vector(-7998,14),
		conv_std_logic_vector(-7999,14),
		conv_std_logic_vector(-8001,14),
		conv_std_logic_vector(-8002,14),
		conv_std_logic_vector(-8003,14),
		conv_std_logic_vector(-8005,14),
		conv_std_logic_vector(-8006,14),
		conv_std_logic_vector(-8007,14),
		conv_std_logic_vector(-8009,14),
		conv_std_logic_vector(-8010,14),
		conv_std_logic_vector(-8011,14),
		conv_std_logic_vector(-8013,14),
		conv_std_logic_vector(-8014,14),
		conv_std_logic_vector(-8015,14),
		conv_std_logic_vector(-8016,14),
		conv_std_logic_vector(-8018,14),
		conv_std_logic_vector(-8019,14),
		conv_std_logic_vector(-8020,14),
		conv_std_logic_vector(-8022,14),
		conv_std_logic_vector(-8023,14),
		conv_std_logic_vector(-8024,14),
		conv_std_logic_vector(-8025,14),
		conv_std_logic_vector(-8027,14),
		conv_std_logic_vector(-8028,14),
		conv_std_logic_vector(-8029,14),
		conv_std_logic_vector(-8030,14),
		conv_std_logic_vector(-8032,14),
		conv_std_logic_vector(-8033,14),
		conv_std_logic_vector(-8034,14),
		conv_std_logic_vector(-8035,14),
		conv_std_logic_vector(-8037,14),
		conv_std_logic_vector(-8038,14),
		conv_std_logic_vector(-8039,14),
		conv_std_logic_vector(-8040,14),
		conv_std_logic_vector(-8041,14),
		conv_std_logic_vector(-8043,14),
		conv_std_logic_vector(-8044,14),
		conv_std_logic_vector(-8045,14),
		conv_std_logic_vector(-8046,14),
		conv_std_logic_vector(-8047,14),
		conv_std_logic_vector(-8048,14),
		conv_std_logic_vector(-8050,14),
		conv_std_logic_vector(-8051,14),
		conv_std_logic_vector(-8052,14),
		conv_std_logic_vector(-8053,14),
		conv_std_logic_vector(-8054,14),
		conv_std_logic_vector(-8055,14),
		conv_std_logic_vector(-8057,14),
		conv_std_logic_vector(-8058,14),
		conv_std_logic_vector(-8059,14),
		conv_std_logic_vector(-8060,14),
		conv_std_logic_vector(-8061,14),
		conv_std_logic_vector(-8062,14),
		conv_std_logic_vector(-8063,14),
		conv_std_logic_vector(-8064,14),
		conv_std_logic_vector(-8065,14),
		conv_std_logic_vector(-8067,14),
		conv_std_logic_vector(-8068,14),
		conv_std_logic_vector(-8069,14),
		conv_std_logic_vector(-8070,14),
		conv_std_logic_vector(-8071,14),
		conv_std_logic_vector(-8072,14),
		conv_std_logic_vector(-8073,14),
		conv_std_logic_vector(-8074,14),
		conv_std_logic_vector(-8075,14),
		conv_std_logic_vector(-8076,14),
		conv_std_logic_vector(-8077,14),
		conv_std_logic_vector(-8078,14),
		conv_std_logic_vector(-8079,14),
		conv_std_logic_vector(-8080,14),
		conv_std_logic_vector(-8081,14),
		conv_std_logic_vector(-8082,14),
		conv_std_logic_vector(-8083,14),
		conv_std_logic_vector(-8084,14),
		conv_std_logic_vector(-8085,14),
		conv_std_logic_vector(-8086,14),
		conv_std_logic_vector(-8087,14),
		conv_std_logic_vector(-8088,14),
		conv_std_logic_vector(-8089,14),
		conv_std_logic_vector(-8090,14),
		conv_std_logic_vector(-8091,14),
		conv_std_logic_vector(-8092,14),
		conv_std_logic_vector(-8093,14),
		conv_std_logic_vector(-8094,14),
		conv_std_logic_vector(-8095,14),
		conv_std_logic_vector(-8096,14),
		conv_std_logic_vector(-8097,14),
		conv_std_logic_vector(-8098,14),
		conv_std_logic_vector(-8099,14),
		conv_std_logic_vector(-8100,14),
		conv_std_logic_vector(-8101,14),
		conv_std_logic_vector(-8102,14),
		conv_std_logic_vector(-8103,14),
		conv_std_logic_vector(-8104,14),
		conv_std_logic_vector(-8105,14),
		conv_std_logic_vector(-8106,14),
		conv_std_logic_vector(-8106,14),
		conv_std_logic_vector(-8107,14),
		conv_std_logic_vector(-8108,14),
		conv_std_logic_vector(-8109,14),
		conv_std_logic_vector(-8110,14),
		conv_std_logic_vector(-8111,14),
		conv_std_logic_vector(-8112,14),
		conv_std_logic_vector(-8113,14),
		conv_std_logic_vector(-8114,14),
		conv_std_logic_vector(-8114,14),
		conv_std_logic_vector(-8115,14),
		conv_std_logic_vector(-8116,14),
		conv_std_logic_vector(-8117,14),
		conv_std_logic_vector(-8118,14),
		conv_std_logic_vector(-8119,14),
		conv_std_logic_vector(-8119,14),
		conv_std_logic_vector(-8120,14),
		conv_std_logic_vector(-8121,14),
		conv_std_logic_vector(-8122,14),
		conv_std_logic_vector(-8123,14),
		conv_std_logic_vector(-8124,14),
		conv_std_logic_vector(-8124,14),
		conv_std_logic_vector(-8125,14),
		conv_std_logic_vector(-8126,14),
		conv_std_logic_vector(-8127,14),
		conv_std_logic_vector(-8128,14),
		conv_std_logic_vector(-8128,14),
		conv_std_logic_vector(-8129,14),
		conv_std_logic_vector(-8130,14),
		conv_std_logic_vector(-8131,14),
		conv_std_logic_vector(-8131,14),
		conv_std_logic_vector(-8132,14),
		conv_std_logic_vector(-8133,14),
		conv_std_logic_vector(-8134,14),
		conv_std_logic_vector(-8134,14),
		conv_std_logic_vector(-8135,14),
		conv_std_logic_vector(-8136,14),
		conv_std_logic_vector(-8137,14),
		conv_std_logic_vector(-8137,14),
		conv_std_logic_vector(-8138,14),
		conv_std_logic_vector(-8139,14),
		conv_std_logic_vector(-8139,14),
		conv_std_logic_vector(-8140,14),
		conv_std_logic_vector(-8141,14),
		conv_std_logic_vector(-8142,14),
		conv_std_logic_vector(-8142,14),
		conv_std_logic_vector(-8143,14),
		conv_std_logic_vector(-8144,14),
		conv_std_logic_vector(-8144,14),
		conv_std_logic_vector(-8145,14),
		conv_std_logic_vector(-8146,14),
		conv_std_logic_vector(-8146,14),
		conv_std_logic_vector(-8147,14),
		conv_std_logic_vector(-8148,14),
		conv_std_logic_vector(-8148,14),
		conv_std_logic_vector(-8149,14),
		conv_std_logic_vector(-8150,14),
		conv_std_logic_vector(-8150,14),
		conv_std_logic_vector(-8151,14),
		conv_std_logic_vector(-8151,14),
		conv_std_logic_vector(-8152,14),
		conv_std_logic_vector(-8153,14),
		conv_std_logic_vector(-8153,14),
		conv_std_logic_vector(-8154,14),
		conv_std_logic_vector(-8154,14),
		conv_std_logic_vector(-8155,14),
		conv_std_logic_vector(-8156,14),
		conv_std_logic_vector(-8156,14),
		conv_std_logic_vector(-8157,14),
		conv_std_logic_vector(-8157,14),
		conv_std_logic_vector(-8158,14),
		conv_std_logic_vector(-8159,14),
		conv_std_logic_vector(-8159,14),
		conv_std_logic_vector(-8160,14),
		conv_std_logic_vector(-8160,14),
		conv_std_logic_vector(-8161,14),
		conv_std_logic_vector(-8161,14),
		conv_std_logic_vector(-8162,14),
		conv_std_logic_vector(-8162,14),
		conv_std_logic_vector(-8163,14),
		conv_std_logic_vector(-8163,14),
		conv_std_logic_vector(-8164,14),
		conv_std_logic_vector(-8164,14),
		conv_std_logic_vector(-8165,14),
		conv_std_logic_vector(-8165,14),
		conv_std_logic_vector(-8166,14),
		conv_std_logic_vector(-8166,14),
		conv_std_logic_vector(-8167,14),
		conv_std_logic_vector(-8167,14),
		conv_std_logic_vector(-8168,14),
		conv_std_logic_vector(-8168,14),
		conv_std_logic_vector(-8169,14),
		conv_std_logic_vector(-8169,14),
		conv_std_logic_vector(-8170,14),
		conv_std_logic_vector(-8170,14),
		conv_std_logic_vector(-8171,14),
		conv_std_logic_vector(-8171,14),
		conv_std_logic_vector(-8172,14),
		conv_std_logic_vector(-8172,14),
		conv_std_logic_vector(-8172,14),
		conv_std_logic_vector(-8173,14),
		conv_std_logic_vector(-8173,14),
		conv_std_logic_vector(-8174,14),
		conv_std_logic_vector(-8174,14),
		conv_std_logic_vector(-8175,14),
		conv_std_logic_vector(-8175,14),
		conv_std_logic_vector(-8175,14),
		conv_std_logic_vector(-8176,14),
		conv_std_logic_vector(-8176,14),
		conv_std_logic_vector(-8176,14),
		conv_std_logic_vector(-8177,14),
		conv_std_logic_vector(-8177,14),
		conv_std_logic_vector(-8178,14),
		conv_std_logic_vector(-8178,14),
		conv_std_logic_vector(-8178,14),
		conv_std_logic_vector(-8179,14),
		conv_std_logic_vector(-8179,14),
		conv_std_logic_vector(-8179,14),
		conv_std_logic_vector(-8180,14),
		conv_std_logic_vector(-8180,14),
		conv_std_logic_vector(-8180,14),
		conv_std_logic_vector(-8181,14),
		conv_std_logic_vector(-8181,14),
		conv_std_logic_vector(-8181,14),
		conv_std_logic_vector(-8182,14),
		conv_std_logic_vector(-8182,14),
		conv_std_logic_vector(-8182,14),
		conv_std_logic_vector(-8183,14),
		conv_std_logic_vector(-8183,14),
		conv_std_logic_vector(-8183,14),
		conv_std_logic_vector(-8183,14),
		conv_std_logic_vector(-8184,14),
		conv_std_logic_vector(-8184,14),
		conv_std_logic_vector(-8184,14),
		conv_std_logic_vector(-8184,14),
		conv_std_logic_vector(-8185,14),
		conv_std_logic_vector(-8185,14),
		conv_std_logic_vector(-8185,14),
		conv_std_logic_vector(-8185,14),
		conv_std_logic_vector(-8186,14),
		conv_std_logic_vector(-8186,14),
		conv_std_logic_vector(-8186,14),
		conv_std_logic_vector(-8186,14),
		conv_std_logic_vector(-8187,14),
		conv_std_logic_vector(-8187,14),
		conv_std_logic_vector(-8187,14),
		conv_std_logic_vector(-8187,14),
		conv_std_logic_vector(-8187,14),
		conv_std_logic_vector(-8188,14),
		conv_std_logic_vector(-8188,14),
		conv_std_logic_vector(-8188,14),
		conv_std_logic_vector(-8188,14),
		conv_std_logic_vector(-8188,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8192,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8191,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8190,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8189,14),
		conv_std_logic_vector(-8188,14),
		conv_std_logic_vector(-8188,14),
		conv_std_logic_vector(-8188,14),
		conv_std_logic_vector(-8188,14),
		conv_std_logic_vector(-8188,14),
		conv_std_logic_vector(-8187,14),
		conv_std_logic_vector(-8187,14),
		conv_std_logic_vector(-8187,14),
		conv_std_logic_vector(-8187,14),
		conv_std_logic_vector(-8187,14),
		conv_std_logic_vector(-8186,14),
		conv_std_logic_vector(-8186,14),
		conv_std_logic_vector(-8186,14),
		conv_std_logic_vector(-8186,14),
		conv_std_logic_vector(-8185,14),
		conv_std_logic_vector(-8185,14),
		conv_std_logic_vector(-8185,14),
		conv_std_logic_vector(-8185,14),
		conv_std_logic_vector(-8184,14),
		conv_std_logic_vector(-8184,14),
		conv_std_logic_vector(-8184,14),
		conv_std_logic_vector(-8184,14),
		conv_std_logic_vector(-8183,14),
		conv_std_logic_vector(-8183,14),
		conv_std_logic_vector(-8183,14),
		conv_std_logic_vector(-8183,14),
		conv_std_logic_vector(-8182,14),
		conv_std_logic_vector(-8182,14),
		conv_std_logic_vector(-8182,14),
		conv_std_logic_vector(-8181,14),
		conv_std_logic_vector(-8181,14),
		conv_std_logic_vector(-8181,14),
		conv_std_logic_vector(-8180,14),
		conv_std_logic_vector(-8180,14),
		conv_std_logic_vector(-8180,14),
		conv_std_logic_vector(-8179,14),
		conv_std_logic_vector(-8179,14),
		conv_std_logic_vector(-8179,14),
		conv_std_logic_vector(-8178,14),
		conv_std_logic_vector(-8178,14),
		conv_std_logic_vector(-8178,14),
		conv_std_logic_vector(-8177,14),
		conv_std_logic_vector(-8177,14),
		conv_std_logic_vector(-8176,14),
		conv_std_logic_vector(-8176,14),
		conv_std_logic_vector(-8176,14),
		conv_std_logic_vector(-8175,14),
		conv_std_logic_vector(-8175,14),
		conv_std_logic_vector(-8175,14),
		conv_std_logic_vector(-8174,14),
		conv_std_logic_vector(-8174,14),
		conv_std_logic_vector(-8173,14),
		conv_std_logic_vector(-8173,14),
		conv_std_logic_vector(-8172,14),
		conv_std_logic_vector(-8172,14),
		conv_std_logic_vector(-8172,14),
		conv_std_logic_vector(-8171,14),
		conv_std_logic_vector(-8171,14),
		conv_std_logic_vector(-8170,14),
		conv_std_logic_vector(-8170,14),
		conv_std_logic_vector(-8169,14),
		conv_std_logic_vector(-8169,14),
		conv_std_logic_vector(-8168,14),
		conv_std_logic_vector(-8168,14),
		conv_std_logic_vector(-8167,14),
		conv_std_logic_vector(-8167,14),
		conv_std_logic_vector(-8166,14),
		conv_std_logic_vector(-8166,14),
		conv_std_logic_vector(-8165,14),
		conv_std_logic_vector(-8165,14),
		conv_std_logic_vector(-8164,14),
		conv_std_logic_vector(-8164,14),
		conv_std_logic_vector(-8163,14),
		conv_std_logic_vector(-8163,14),
		conv_std_logic_vector(-8162,14),
		conv_std_logic_vector(-8162,14),
		conv_std_logic_vector(-8161,14),
		conv_std_logic_vector(-8161,14),
		conv_std_logic_vector(-8160,14),
		conv_std_logic_vector(-8160,14),
		conv_std_logic_vector(-8159,14),
		conv_std_logic_vector(-8159,14),
		conv_std_logic_vector(-8158,14),
		conv_std_logic_vector(-8157,14),
		conv_std_logic_vector(-8157,14),
		conv_std_logic_vector(-8156,14),
		conv_std_logic_vector(-8156,14),
		conv_std_logic_vector(-8155,14),
		conv_std_logic_vector(-8154,14),
		conv_std_logic_vector(-8154,14),
		conv_std_logic_vector(-8153,14),
		conv_std_logic_vector(-8153,14),
		conv_std_logic_vector(-8152,14),
		conv_std_logic_vector(-8151,14),
		conv_std_logic_vector(-8151,14),
		conv_std_logic_vector(-8150,14),
		conv_std_logic_vector(-8150,14),
		conv_std_logic_vector(-8149,14),
		conv_std_logic_vector(-8148,14),
		conv_std_logic_vector(-8148,14),
		conv_std_logic_vector(-8147,14),
		conv_std_logic_vector(-8146,14),
		conv_std_logic_vector(-8146,14),
		conv_std_logic_vector(-8145,14),
		conv_std_logic_vector(-8144,14),
		conv_std_logic_vector(-8144,14),
		conv_std_logic_vector(-8143,14),
		conv_std_logic_vector(-8142,14),
		conv_std_logic_vector(-8142,14),
		conv_std_logic_vector(-8141,14),
		conv_std_logic_vector(-8140,14),
		conv_std_logic_vector(-8139,14),
		conv_std_logic_vector(-8139,14),
		conv_std_logic_vector(-8138,14),
		conv_std_logic_vector(-8137,14),
		conv_std_logic_vector(-8137,14),
		conv_std_logic_vector(-8136,14),
		conv_std_logic_vector(-8135,14),
		conv_std_logic_vector(-8134,14),
		conv_std_logic_vector(-8134,14),
		conv_std_logic_vector(-8133,14),
		conv_std_logic_vector(-8132,14),
		conv_std_logic_vector(-8131,14),
		conv_std_logic_vector(-8131,14),
		conv_std_logic_vector(-8130,14),
		conv_std_logic_vector(-8129,14),
		conv_std_logic_vector(-8128,14),
		conv_std_logic_vector(-8128,14),
		conv_std_logic_vector(-8127,14),
		conv_std_logic_vector(-8126,14),
		conv_std_logic_vector(-8125,14),
		conv_std_logic_vector(-8124,14),
		conv_std_logic_vector(-8124,14),
		conv_std_logic_vector(-8123,14),
		conv_std_logic_vector(-8122,14),
		conv_std_logic_vector(-8121,14),
		conv_std_logic_vector(-8120,14),
		conv_std_logic_vector(-8119,14),
		conv_std_logic_vector(-8119,14),
		conv_std_logic_vector(-8118,14),
		conv_std_logic_vector(-8117,14),
		conv_std_logic_vector(-8116,14),
		conv_std_logic_vector(-8115,14),
		conv_std_logic_vector(-8114,14),
		conv_std_logic_vector(-8114,14),
		conv_std_logic_vector(-8113,14),
		conv_std_logic_vector(-8112,14),
		conv_std_logic_vector(-8111,14),
		conv_std_logic_vector(-8110,14),
		conv_std_logic_vector(-8109,14),
		conv_std_logic_vector(-8108,14),
		conv_std_logic_vector(-8107,14),
		conv_std_logic_vector(-8106,14),
		conv_std_logic_vector(-8106,14),
		conv_std_logic_vector(-8105,14),
		conv_std_logic_vector(-8104,14),
		conv_std_logic_vector(-8103,14),
		conv_std_logic_vector(-8102,14),
		conv_std_logic_vector(-8101,14),
		conv_std_logic_vector(-8100,14),
		conv_std_logic_vector(-8099,14),
		conv_std_logic_vector(-8098,14),
		conv_std_logic_vector(-8097,14),
		conv_std_logic_vector(-8096,14),
		conv_std_logic_vector(-8095,14),
		conv_std_logic_vector(-8094,14),
		conv_std_logic_vector(-8093,14),
		conv_std_logic_vector(-8092,14),
		conv_std_logic_vector(-8091,14),
		conv_std_logic_vector(-8090,14),
		conv_std_logic_vector(-8089,14),
		conv_std_logic_vector(-8088,14),
		conv_std_logic_vector(-8087,14),
		conv_std_logic_vector(-8086,14),
		conv_std_logic_vector(-8085,14),
		conv_std_logic_vector(-8084,14),
		conv_std_logic_vector(-8083,14),
		conv_std_logic_vector(-8082,14),
		conv_std_logic_vector(-8081,14),
		conv_std_logic_vector(-8080,14),
		conv_std_logic_vector(-8079,14),
		conv_std_logic_vector(-8078,14),
		conv_std_logic_vector(-8077,14),
		conv_std_logic_vector(-8076,14),
		conv_std_logic_vector(-8075,14),
		conv_std_logic_vector(-8074,14),
		conv_std_logic_vector(-8073,14),
		conv_std_logic_vector(-8072,14),
		conv_std_logic_vector(-8071,14),
		conv_std_logic_vector(-8070,14),
		conv_std_logic_vector(-8069,14),
		conv_std_logic_vector(-8068,14),
		conv_std_logic_vector(-8067,14),
		conv_std_logic_vector(-8065,14),
		conv_std_logic_vector(-8064,14),
		conv_std_logic_vector(-8063,14),
		conv_std_logic_vector(-8062,14),
		conv_std_logic_vector(-8061,14),
		conv_std_logic_vector(-8060,14),
		conv_std_logic_vector(-8059,14),
		conv_std_logic_vector(-8058,14),
		conv_std_logic_vector(-8057,14),
		conv_std_logic_vector(-8055,14),
		conv_std_logic_vector(-8054,14),
		conv_std_logic_vector(-8053,14),
		conv_std_logic_vector(-8052,14),
		conv_std_logic_vector(-8051,14),
		conv_std_logic_vector(-8050,14),
		conv_std_logic_vector(-8048,14),
		conv_std_logic_vector(-8047,14),
		conv_std_logic_vector(-8046,14),
		conv_std_logic_vector(-8045,14),
		conv_std_logic_vector(-8044,14),
		conv_std_logic_vector(-8043,14),
		conv_std_logic_vector(-8041,14),
		conv_std_logic_vector(-8040,14),
		conv_std_logic_vector(-8039,14),
		conv_std_logic_vector(-8038,14),
		conv_std_logic_vector(-8037,14),
		conv_std_logic_vector(-8035,14),
		conv_std_logic_vector(-8034,14),
		conv_std_logic_vector(-8033,14),
		conv_std_logic_vector(-8032,14),
		conv_std_logic_vector(-8030,14),
		conv_std_logic_vector(-8029,14),
		conv_std_logic_vector(-8028,14),
		conv_std_logic_vector(-8027,14),
		conv_std_logic_vector(-8025,14),
		conv_std_logic_vector(-8024,14),
		conv_std_logic_vector(-8023,14),
		conv_std_logic_vector(-8022,14),
		conv_std_logic_vector(-8020,14),
		conv_std_logic_vector(-8019,14),
		conv_std_logic_vector(-8018,14),
		conv_std_logic_vector(-8016,14),
		conv_std_logic_vector(-8015,14),
		conv_std_logic_vector(-8014,14),
		conv_std_logic_vector(-8013,14),
		conv_std_logic_vector(-8011,14),
		conv_std_logic_vector(-8010,14),
		conv_std_logic_vector(-8009,14),
		conv_std_logic_vector(-8007,14),
		conv_std_logic_vector(-8006,14),
		conv_std_logic_vector(-8005,14),
		conv_std_logic_vector(-8003,14),
		conv_std_logic_vector(-8002,14),
		conv_std_logic_vector(-8001,14),
		conv_std_logic_vector(-7999,14),
		conv_std_logic_vector(-7998,14),
		conv_std_logic_vector(-7997,14),
		conv_std_logic_vector(-7995,14),
		conv_std_logic_vector(-7994,14),
		conv_std_logic_vector(-7992,14),
		conv_std_logic_vector(-7991,14),
		conv_std_logic_vector(-7990,14),
		conv_std_logic_vector(-7988,14),
		conv_std_logic_vector(-7987,14),
		conv_std_logic_vector(-7986,14),
		conv_std_logic_vector(-7984,14),
		conv_std_logic_vector(-7983,14),
		conv_std_logic_vector(-7981,14),
		conv_std_logic_vector(-7980,14),
		conv_std_logic_vector(-7978,14),
		conv_std_logic_vector(-7977,14),
		conv_std_logic_vector(-7976,14),
		conv_std_logic_vector(-7974,14),
		conv_std_logic_vector(-7973,14),
		conv_std_logic_vector(-7971,14),
		conv_std_logic_vector(-7970,14),
		conv_std_logic_vector(-7968,14),
		conv_std_logic_vector(-7967,14),
		conv_std_logic_vector(-7965,14),
		conv_std_logic_vector(-7964,14),
		conv_std_logic_vector(-7963,14),
		conv_std_logic_vector(-7961,14),
		conv_std_logic_vector(-7960,14),
		conv_std_logic_vector(-7958,14),
		conv_std_logic_vector(-7957,14),
		conv_std_logic_vector(-7955,14),
		conv_std_logic_vector(-7954,14),
		conv_std_logic_vector(-7952,14),
		conv_std_logic_vector(-7951,14),
		conv_std_logic_vector(-7949,14),
		conv_std_logic_vector(-7948,14),
		conv_std_logic_vector(-7946,14),
		conv_std_logic_vector(-7944,14),
		conv_std_logic_vector(-7943,14),
		conv_std_logic_vector(-7941,14),
		conv_std_logic_vector(-7940,14),
		conv_std_logic_vector(-7938,14),
		conv_std_logic_vector(-7937,14),
		conv_std_logic_vector(-7935,14),
		conv_std_logic_vector(-7934,14),
		conv_std_logic_vector(-7932,14),
		conv_std_logic_vector(-7930,14),
		conv_std_logic_vector(-7929,14),
		conv_std_logic_vector(-7927,14),
		conv_std_logic_vector(-7926,14),
		conv_std_logic_vector(-7924,14),
		conv_std_logic_vector(-7923,14),
		conv_std_logic_vector(-7921,14),
		conv_std_logic_vector(-7919,14),
		conv_std_logic_vector(-7918,14),
		conv_std_logic_vector(-7916,14),
		conv_std_logic_vector(-7915,14),
		conv_std_logic_vector(-7913,14),
		conv_std_logic_vector(-7911,14),
		conv_std_logic_vector(-7910,14),
		conv_std_logic_vector(-7908,14),
		conv_std_logic_vector(-7906,14),
		conv_std_logic_vector(-7905,14),
		conv_std_logic_vector(-7903,14),
		conv_std_logic_vector(-7901,14),
		conv_std_logic_vector(-7900,14),
		conv_std_logic_vector(-7898,14),
		conv_std_logic_vector(-7896,14),
		conv_std_logic_vector(-7895,14),
		conv_std_logic_vector(-7893,14),
		conv_std_logic_vector(-7891,14),
		conv_std_logic_vector(-7890,14),
		conv_std_logic_vector(-7888,14),
		conv_std_logic_vector(-7886,14),
		conv_std_logic_vector(-7885,14),
		conv_std_logic_vector(-7883,14),
		conv_std_logic_vector(-7881,14),
		conv_std_logic_vector(-7879,14),
		conv_std_logic_vector(-7878,14),
		conv_std_logic_vector(-7876,14),
		conv_std_logic_vector(-7874,14),
		conv_std_logic_vector(-7873,14),
		conv_std_logic_vector(-7871,14),
		conv_std_logic_vector(-7869,14),
		conv_std_logic_vector(-7867,14),
		conv_std_logic_vector(-7866,14),
		conv_std_logic_vector(-7864,14),
		conv_std_logic_vector(-7862,14),
		conv_std_logic_vector(-7860,14),
		conv_std_logic_vector(-7859,14),
		conv_std_logic_vector(-7857,14),
		conv_std_logic_vector(-7855,14),
		conv_std_logic_vector(-7853,14),
		conv_std_logic_vector(-7851,14),
		conv_std_logic_vector(-7850,14),
		conv_std_logic_vector(-7848,14),
		conv_std_logic_vector(-7846,14),
		conv_std_logic_vector(-7844,14),
		conv_std_logic_vector(-7842,14),
		conv_std_logic_vector(-7841,14),
		conv_std_logic_vector(-7839,14),
		conv_std_logic_vector(-7837,14),
		conv_std_logic_vector(-7835,14),
		conv_std_logic_vector(-7833,14),
		conv_std_logic_vector(-7831,14),
		conv_std_logic_vector(-7830,14),
		conv_std_logic_vector(-7828,14),
		conv_std_logic_vector(-7826,14),
		conv_std_logic_vector(-7824,14),
		conv_std_logic_vector(-7822,14),
		conv_std_logic_vector(-7820,14),
		conv_std_logic_vector(-7818,14),
		conv_std_logic_vector(-7817,14),
		conv_std_logic_vector(-7815,14),
		conv_std_logic_vector(-7813,14),
		conv_std_logic_vector(-7811,14),
		conv_std_logic_vector(-7809,14),
		conv_std_logic_vector(-7807,14),
		conv_std_logic_vector(-7805,14),
		conv_std_logic_vector(-7803,14),
		conv_std_logic_vector(-7801,14),
		conv_std_logic_vector(-7799,14),
		conv_std_logic_vector(-7798,14),
		conv_std_logic_vector(-7796,14),
		conv_std_logic_vector(-7794,14),
		conv_std_logic_vector(-7792,14),
		conv_std_logic_vector(-7790,14),
		conv_std_logic_vector(-7788,14),
		conv_std_logic_vector(-7786,14),
		conv_std_logic_vector(-7784,14),
		conv_std_logic_vector(-7782,14),
		conv_std_logic_vector(-7780,14),
		conv_std_logic_vector(-7778,14),
		conv_std_logic_vector(-7776,14),
		conv_std_logic_vector(-7774,14),
		conv_std_logic_vector(-7772,14),
		conv_std_logic_vector(-7770,14),
		conv_std_logic_vector(-7768,14),
		conv_std_logic_vector(-7766,14),
		conv_std_logic_vector(-7764,14),
		conv_std_logic_vector(-7762,14),
		conv_std_logic_vector(-7760,14),
		conv_std_logic_vector(-7758,14),
		conv_std_logic_vector(-7756,14),
		conv_std_logic_vector(-7754,14),
		conv_std_logic_vector(-7752,14),
		conv_std_logic_vector(-7750,14),
		conv_std_logic_vector(-7748,14),
		conv_std_logic_vector(-7746,14),
		conv_std_logic_vector(-7744,14),
		conv_std_logic_vector(-7742,14),
		conv_std_logic_vector(-7740,14),
		conv_std_logic_vector(-7738,14),
		conv_std_logic_vector(-7736,14),
		conv_std_logic_vector(-7734,14),
		conv_std_logic_vector(-7731,14),
		conv_std_logic_vector(-7729,14),
		conv_std_logic_vector(-7727,14),
		conv_std_logic_vector(-7725,14),
		conv_std_logic_vector(-7723,14),
		conv_std_logic_vector(-7721,14),
		conv_std_logic_vector(-7719,14),
		conv_std_logic_vector(-7717,14),
		conv_std_logic_vector(-7715,14),
		conv_std_logic_vector(-7713,14),
		conv_std_logic_vector(-7711,14),
		conv_std_logic_vector(-7708,14),
		conv_std_logic_vector(-7706,14),
		conv_std_logic_vector(-7704,14),
		conv_std_logic_vector(-7702,14),
		conv_std_logic_vector(-7700,14),
		conv_std_logic_vector(-7698,14),
		conv_std_logic_vector(-7696,14),
		conv_std_logic_vector(-7693,14),
		conv_std_logic_vector(-7691,14),
		conv_std_logic_vector(-7689,14),
		conv_std_logic_vector(-7687,14),
		conv_std_logic_vector(-7685,14),
		conv_std_logic_vector(-7683,14),
		conv_std_logic_vector(-7680,14),
		conv_std_logic_vector(-7678,14),
		conv_std_logic_vector(-7676,14),
		conv_std_logic_vector(-7674,14),
		conv_std_logic_vector(-7672,14),
		conv_std_logic_vector(-7669,14),
		conv_std_logic_vector(-7667,14),
		conv_std_logic_vector(-7665,14),
		conv_std_logic_vector(-7663,14),
		conv_std_logic_vector(-7661,14),
		conv_std_logic_vector(-7658,14),
		conv_std_logic_vector(-7656,14),
		conv_std_logic_vector(-7654,14),
		conv_std_logic_vector(-7652,14),
		conv_std_logic_vector(-7649,14),
		conv_std_logic_vector(-7647,14),
		conv_std_logic_vector(-7645,14),
		conv_std_logic_vector(-7643,14),
		conv_std_logic_vector(-7640,14),
		conv_std_logic_vector(-7638,14),
		conv_std_logic_vector(-7636,14),
		conv_std_logic_vector(-7633,14),
		conv_std_logic_vector(-7631,14),
		conv_std_logic_vector(-7629,14),
		conv_std_logic_vector(-7627,14),
		conv_std_logic_vector(-7624,14),
		conv_std_logic_vector(-7622,14),
		conv_std_logic_vector(-7620,14),
		conv_std_logic_vector(-7617,14),
		conv_std_logic_vector(-7615,14),
		conv_std_logic_vector(-7613,14),
		conv_std_logic_vector(-7610,14),
		conv_std_logic_vector(-7608,14),
		conv_std_logic_vector(-7606,14),
		conv_std_logic_vector(-7603,14),
		conv_std_logic_vector(-7601,14),
		conv_std_logic_vector(-7599,14),
		conv_std_logic_vector(-7596,14),
		conv_std_logic_vector(-7594,14),
		conv_std_logic_vector(-7592,14),
		conv_std_logic_vector(-7589,14),
		conv_std_logic_vector(-7587,14),
		conv_std_logic_vector(-7585,14),
		conv_std_logic_vector(-7582,14),
		conv_std_logic_vector(-7580,14),
		conv_std_logic_vector(-7578,14),
		conv_std_logic_vector(-7575,14),
		conv_std_logic_vector(-7573,14),
		conv_std_logic_vector(-7570,14),
		conv_std_logic_vector(-7568,14),
		conv_std_logic_vector(-7566,14),
		conv_std_logic_vector(-7563,14),
		conv_std_logic_vector(-7561,14),
		conv_std_logic_vector(-7558,14),
		conv_std_logic_vector(-7556,14),
		conv_std_logic_vector(-7553,14),
		conv_std_logic_vector(-7551,14),
		conv_std_logic_vector(-7549,14),
		conv_std_logic_vector(-7546,14),
		conv_std_logic_vector(-7544,14),
		conv_std_logic_vector(-7541,14),
		conv_std_logic_vector(-7539,14),
		conv_std_logic_vector(-7536,14),
		conv_std_logic_vector(-7534,14),
		conv_std_logic_vector(-7531,14),
		conv_std_logic_vector(-7529,14),
		conv_std_logic_vector(-7526,14),
		conv_std_logic_vector(-7524,14),
		conv_std_logic_vector(-7521,14),
		conv_std_logic_vector(-7519,14),
		conv_std_logic_vector(-7516,14),
		conv_std_logic_vector(-7514,14),
		conv_std_logic_vector(-7511,14),
		conv_std_logic_vector(-7509,14),
		conv_std_logic_vector(-7506,14),
		conv_std_logic_vector(-7504,14),
		conv_std_logic_vector(-7501,14),
		conv_std_logic_vector(-7499,14),
		conv_std_logic_vector(-7496,14),
		conv_std_logic_vector(-7494,14),
		conv_std_logic_vector(-7491,14),
		conv_std_logic_vector(-7489,14),
		conv_std_logic_vector(-7486,14),
		conv_std_logic_vector(-7484,14),
		conv_std_logic_vector(-7481,14),
		conv_std_logic_vector(-7478,14),
		conv_std_logic_vector(-7476,14),
		conv_std_logic_vector(-7473,14),
		conv_std_logic_vector(-7471,14),
		conv_std_logic_vector(-7468,14),
		conv_std_logic_vector(-7466,14),
		conv_std_logic_vector(-7463,14),
		conv_std_logic_vector(-7460,14),
		conv_std_logic_vector(-7458,14),
		conv_std_logic_vector(-7455,14),
		conv_std_logic_vector(-7453,14),
		conv_std_logic_vector(-7450,14),
		conv_std_logic_vector(-7447,14),
		conv_std_logic_vector(-7445,14),
		conv_std_logic_vector(-7442,14),
		conv_std_logic_vector(-7440,14),
		conv_std_logic_vector(-7437,14),
		conv_std_logic_vector(-7434,14),
		conv_std_logic_vector(-7432,14),
		conv_std_logic_vector(-7429,14),
		conv_std_logic_vector(-7426,14),
		conv_std_logic_vector(-7424,14),
		conv_std_logic_vector(-7421,14),
		conv_std_logic_vector(-7418,14),
		conv_std_logic_vector(-7416,14),
		conv_std_logic_vector(-7413,14),
		conv_std_logic_vector(-7410,14),
		conv_std_logic_vector(-7408,14),
		conv_std_logic_vector(-7405,14),
		conv_std_logic_vector(-7402,14),
		conv_std_logic_vector(-7400,14),
		conv_std_logic_vector(-7397,14),
		conv_std_logic_vector(-7394,14),
		conv_std_logic_vector(-7391,14),
		conv_std_logic_vector(-7389,14),
		conv_std_logic_vector(-7386,14),
		conv_std_logic_vector(-7383,14),
		conv_std_logic_vector(-7381,14),
		conv_std_logic_vector(-7378,14),
		conv_std_logic_vector(-7375,14),
		conv_std_logic_vector(-7372,14),
		conv_std_logic_vector(-7370,14),
		conv_std_logic_vector(-7367,14),
		conv_std_logic_vector(-7364,14),
		conv_std_logic_vector(-7361,14),
		conv_std_logic_vector(-7359,14),
		conv_std_logic_vector(-7356,14),
		conv_std_logic_vector(-7353,14),
		conv_std_logic_vector(-7350,14),
		conv_std_logic_vector(-7348,14),
		conv_std_logic_vector(-7345,14),
		conv_std_logic_vector(-7342,14),
		conv_std_logic_vector(-7339,14),
		conv_std_logic_vector(-7336,14),
		conv_std_logic_vector(-7334,14),
		conv_std_logic_vector(-7331,14),
		conv_std_logic_vector(-7328,14),
		conv_std_logic_vector(-7325,14),
		conv_std_logic_vector(-7322,14),
		conv_std_logic_vector(-7320,14),
		conv_std_logic_vector(-7317,14),
		conv_std_logic_vector(-7314,14),
		conv_std_logic_vector(-7311,14),
		conv_std_logic_vector(-7308,14),
		conv_std_logic_vector(-7305,14),
		conv_std_logic_vector(-7303,14),
		conv_std_logic_vector(-7300,14),
		conv_std_logic_vector(-7297,14),
		conv_std_logic_vector(-7294,14),
		conv_std_logic_vector(-7291,14),
		conv_std_logic_vector(-7288,14),
		conv_std_logic_vector(-7285,14),
		conv_std_logic_vector(-7283,14),
		conv_std_logic_vector(-7280,14),
		conv_std_logic_vector(-7277,14),
		conv_std_logic_vector(-7274,14),
		conv_std_logic_vector(-7271,14),
		conv_std_logic_vector(-7268,14),
		conv_std_logic_vector(-7265,14),
		conv_std_logic_vector(-7262,14),
		conv_std_logic_vector(-7259,14),
		conv_std_logic_vector(-7257,14),
		conv_std_logic_vector(-7254,14),
		conv_std_logic_vector(-7251,14),
		conv_std_logic_vector(-7248,14),
		conv_std_logic_vector(-7245,14),
		conv_std_logic_vector(-7242,14),
		conv_std_logic_vector(-7239,14),
		conv_std_logic_vector(-7236,14),
		conv_std_logic_vector(-7233,14),
		conv_std_logic_vector(-7230,14),
		conv_std_logic_vector(-7227,14),
		conv_std_logic_vector(-7224,14),
		conv_std_logic_vector(-7221,14),
		conv_std_logic_vector(-7218,14),
		conv_std_logic_vector(-7215,14),
		conv_std_logic_vector(-7212,14),
		conv_std_logic_vector(-7209,14),
		conv_std_logic_vector(-7206,14),
		conv_std_logic_vector(-7203,14),
		conv_std_logic_vector(-7200,14),
		conv_std_logic_vector(-7197,14),
		conv_std_logic_vector(-7194,14),
		conv_std_logic_vector(-7191,14),
		conv_std_logic_vector(-7188,14),
		conv_std_logic_vector(-7185,14),
		conv_std_logic_vector(-7182,14),
		conv_std_logic_vector(-7179,14),
		conv_std_logic_vector(-7176,14),
		conv_std_logic_vector(-7173,14),
		conv_std_logic_vector(-7170,14),
		conv_std_logic_vector(-7167,14),
		conv_std_logic_vector(-7164,14),
		conv_std_logic_vector(-7161,14),
		conv_std_logic_vector(-7158,14),
		conv_std_logic_vector(-7155,14),
		conv_std_logic_vector(-7152,14),
		conv_std_logic_vector(-7149,14),
		conv_std_logic_vector(-7146,14),
		conv_std_logic_vector(-7143,14),
		conv_std_logic_vector(-7140,14),
		conv_std_logic_vector(-7137,14),
		conv_std_logic_vector(-7133,14),
		conv_std_logic_vector(-7130,14),
		conv_std_logic_vector(-7127,14),
		conv_std_logic_vector(-7124,14),
		conv_std_logic_vector(-7121,14),
		conv_std_logic_vector(-7118,14),
		conv_std_logic_vector(-7115,14),
		conv_std_logic_vector(-7112,14),
		conv_std_logic_vector(-7109,14),
		conv_std_logic_vector(-7105,14),
		conv_std_logic_vector(-7102,14),
		conv_std_logic_vector(-7099,14),
		conv_std_logic_vector(-7096,14),
		conv_std_logic_vector(-7093,14),
		conv_std_logic_vector(-7090,14),
		conv_std_logic_vector(-7087,14),
		conv_std_logic_vector(-7083,14),
		conv_std_logic_vector(-7080,14),
		conv_std_logic_vector(-7077,14),
		conv_std_logic_vector(-7074,14),
		conv_std_logic_vector(-7071,14),
		conv_std_logic_vector(-7068,14),
		conv_std_logic_vector(-7064,14),
		conv_std_logic_vector(-7061,14),
		conv_std_logic_vector(-7058,14),
		conv_std_logic_vector(-7055,14),
		conv_std_logic_vector(-7052,14),
		conv_std_logic_vector(-7049,14),
		conv_std_logic_vector(-7045,14),
		conv_std_logic_vector(-7042,14),
		conv_std_logic_vector(-7039,14),
		conv_std_logic_vector(-7036,14),
		conv_std_logic_vector(-7032,14),
		conv_std_logic_vector(-7029,14),
		conv_std_logic_vector(-7026,14),
		conv_std_logic_vector(-7023,14),
		conv_std_logic_vector(-7020,14),
		conv_std_logic_vector(-7016,14),
		conv_std_logic_vector(-7013,14),
		conv_std_logic_vector(-7010,14),
		conv_std_logic_vector(-7007,14),
		conv_std_logic_vector(-7003,14),
		conv_std_logic_vector(-7000,14),
		conv_std_logic_vector(-6997,14),
		conv_std_logic_vector(-6994,14),
		conv_std_logic_vector(-6990,14),
		conv_std_logic_vector(-6987,14),
		conv_std_logic_vector(-6984,14),
		conv_std_logic_vector(-6980,14),
		conv_std_logic_vector(-6977,14),
		conv_std_logic_vector(-6974,14),
		conv_std_logic_vector(-6971,14),
		conv_std_logic_vector(-6967,14),
		conv_std_logic_vector(-6964,14),
		conv_std_logic_vector(-6961,14),
		conv_std_logic_vector(-6957,14),
		conv_std_logic_vector(-6954,14),
		conv_std_logic_vector(-6951,14),
		conv_std_logic_vector(-6947,14),
		conv_std_logic_vector(-6944,14),
		conv_std_logic_vector(-6941,14),
		conv_std_logic_vector(-6937,14),
		conv_std_logic_vector(-6934,14),
		conv_std_logic_vector(-6931,14),
		conv_std_logic_vector(-6927,14),
		conv_std_logic_vector(-6924,14),
		conv_std_logic_vector(-6921,14),
		conv_std_logic_vector(-6917,14),
		conv_std_logic_vector(-6914,14),
		conv_std_logic_vector(-6910,14),
		conv_std_logic_vector(-6907,14),
		conv_std_logic_vector(-6904,14),
		conv_std_logic_vector(-6900,14),
		conv_std_logic_vector(-6897,14),
		conv_std_logic_vector(-6894,14),
		conv_std_logic_vector(-6890,14),
		conv_std_logic_vector(-6887,14),
		conv_std_logic_vector(-6883,14),
		conv_std_logic_vector(-6880,14),
		conv_std_logic_vector(-6876,14),
		conv_std_logic_vector(-6873,14),
		conv_std_logic_vector(-6870,14),
		conv_std_logic_vector(-6866,14),
		conv_std_logic_vector(-6863,14),
		conv_std_logic_vector(-6859,14),
		conv_std_logic_vector(-6856,14),
		conv_std_logic_vector(-6852,14),
		conv_std_logic_vector(-6849,14),
		conv_std_logic_vector(-6846,14),
		conv_std_logic_vector(-6842,14),
		conv_std_logic_vector(-6839,14),
		conv_std_logic_vector(-6835,14),
		conv_std_logic_vector(-6832,14),
		conv_std_logic_vector(-6828,14),
		conv_std_logic_vector(-6825,14),
		conv_std_logic_vector(-6821,14),
		conv_std_logic_vector(-6818,14),
		conv_std_logic_vector(-6814,14),
		conv_std_logic_vector(-6811,14),
		conv_std_logic_vector(-6807,14),
		conv_std_logic_vector(-6804,14),
		conv_std_logic_vector(-6800,14),
		conv_std_logic_vector(-6797,14),
		conv_std_logic_vector(-6793,14),
		conv_std_logic_vector(-6790,14),
		conv_std_logic_vector(-6786,14),
		conv_std_logic_vector(-6783,14),
		conv_std_logic_vector(-6779,14),
		conv_std_logic_vector(-6776,14),
		conv_std_logic_vector(-6772,14),
		conv_std_logic_vector(-6769,14),
		conv_std_logic_vector(-6765,14),
		conv_std_logic_vector(-6762,14),
		conv_std_logic_vector(-6758,14),
		conv_std_logic_vector(-6755,14),
		conv_std_logic_vector(-6751,14),
		conv_std_logic_vector(-6747,14),
		conv_std_logic_vector(-6744,14),
		conv_std_logic_vector(-6740,14),
		conv_std_logic_vector(-6737,14),
		conv_std_logic_vector(-6733,14),
		conv_std_logic_vector(-6730,14),
		conv_std_logic_vector(-6726,14),
		conv_std_logic_vector(-6722,14),
		conv_std_logic_vector(-6719,14),
		conv_std_logic_vector(-6715,14),
		conv_std_logic_vector(-6712,14),
		conv_std_logic_vector(-6708,14),
		conv_std_logic_vector(-6704,14),
		conv_std_logic_vector(-6701,14),
		conv_std_logic_vector(-6697,14),
		conv_std_logic_vector(-6694,14),
		conv_std_logic_vector(-6690,14),
		conv_std_logic_vector(-6686,14),
		conv_std_logic_vector(-6683,14),
		conv_std_logic_vector(-6679,14),
		conv_std_logic_vector(-6675,14),
		conv_std_logic_vector(-6672,14),
		conv_std_logic_vector(-6668,14),
		conv_std_logic_vector(-6664,14),
		conv_std_logic_vector(-6661,14),
		conv_std_logic_vector(-6657,14),
		conv_std_logic_vector(-6653,14),
		conv_std_logic_vector(-6650,14),
		conv_std_logic_vector(-6646,14),
		conv_std_logic_vector(-6642,14),
		conv_std_logic_vector(-6639,14),
		conv_std_logic_vector(-6635,14),
		conv_std_logic_vector(-6631,14),
		conv_std_logic_vector(-6628,14),
		conv_std_logic_vector(-6624,14),
		conv_std_logic_vector(-6620,14),
		conv_std_logic_vector(-6617,14),
		conv_std_logic_vector(-6613,14),
		conv_std_logic_vector(-6609,14),
		conv_std_logic_vector(-6605,14),
		conv_std_logic_vector(-6602,14),
		conv_std_logic_vector(-6598,14),
		conv_std_logic_vector(-6594,14),
		conv_std_logic_vector(-6591,14),
		conv_std_logic_vector(-6587,14),
		conv_std_logic_vector(-6583,14),
		conv_std_logic_vector(-6579,14),
		conv_std_logic_vector(-6576,14),
		conv_std_logic_vector(-6572,14),
		conv_std_logic_vector(-6568,14),
		conv_std_logic_vector(-6564,14),
		conv_std_logic_vector(-6561,14),
		conv_std_logic_vector(-6557,14),
		conv_std_logic_vector(-6553,14),
		conv_std_logic_vector(-6549,14),
		conv_std_logic_vector(-6546,14),
		conv_std_logic_vector(-6542,14),
		conv_std_logic_vector(-6538,14),
		conv_std_logic_vector(-6534,14),
		conv_std_logic_vector(-6530,14),
		conv_std_logic_vector(-6527,14),
		conv_std_logic_vector(-6523,14),
		conv_std_logic_vector(-6519,14),
		conv_std_logic_vector(-6515,14),
		conv_std_logic_vector(-6511,14),
		conv_std_logic_vector(-6508,14),
		conv_std_logic_vector(-6504,14),
		conv_std_logic_vector(-6500,14),
		conv_std_logic_vector(-6496,14),
		conv_std_logic_vector(-6492,14),
		conv_std_logic_vector(-6488,14),
		conv_std_logic_vector(-6485,14),
		conv_std_logic_vector(-6481,14),
		conv_std_logic_vector(-6477,14),
		conv_std_logic_vector(-6473,14),
		conv_std_logic_vector(-6469,14),
		conv_std_logic_vector(-6465,14),
		conv_std_logic_vector(-6461,14),
		conv_std_logic_vector(-6458,14),
		conv_std_logic_vector(-6454,14),
		conv_std_logic_vector(-6450,14),
		conv_std_logic_vector(-6446,14),
		conv_std_logic_vector(-6442,14),
		conv_std_logic_vector(-6438,14),
		conv_std_logic_vector(-6434,14),
		conv_std_logic_vector(-6430,14),
		conv_std_logic_vector(-6427,14),
		conv_std_logic_vector(-6423,14),
		conv_std_logic_vector(-6419,14),
		conv_std_logic_vector(-6415,14),
		conv_std_logic_vector(-6411,14),
		conv_std_logic_vector(-6407,14),
		conv_std_logic_vector(-6403,14),
		conv_std_logic_vector(-6399,14),
		conv_std_logic_vector(-6395,14),
		conv_std_logic_vector(-6391,14),
		conv_std_logic_vector(-6387,14),
		conv_std_logic_vector(-6384,14),
		conv_std_logic_vector(-6380,14),
		conv_std_logic_vector(-6376,14),
		conv_std_logic_vector(-6372,14),
		conv_std_logic_vector(-6368,14),
		conv_std_logic_vector(-6364,14),
		conv_std_logic_vector(-6360,14),
		conv_std_logic_vector(-6356,14),
		conv_std_logic_vector(-6352,14),
		conv_std_logic_vector(-6348,14),
		conv_std_logic_vector(-6344,14),
		conv_std_logic_vector(-6340,14),
		conv_std_logic_vector(-6336,14),
		conv_std_logic_vector(-6332,14),
		conv_std_logic_vector(-6328,14),
		conv_std_logic_vector(-6324,14),
		conv_std_logic_vector(-6320,14),
		conv_std_logic_vector(-6316,14),
		conv_std_logic_vector(-6312,14),
		conv_std_logic_vector(-6308,14),
		conv_std_logic_vector(-6304,14),
		conv_std_logic_vector(-6300,14),
		conv_std_logic_vector(-6296,14),
		conv_std_logic_vector(-6292,14),
		conv_std_logic_vector(-6288,14),
		conv_std_logic_vector(-6284,14),
		conv_std_logic_vector(-6280,14),
		conv_std_logic_vector(-6276,14),
		conv_std_logic_vector(-6272,14),
		conv_std_logic_vector(-6268,14),
		conv_std_logic_vector(-6264,14),
		conv_std_logic_vector(-6260,14),
		conv_std_logic_vector(-6256,14),
		conv_std_logic_vector(-6252,14),
		conv_std_logic_vector(-6247,14),
		conv_std_logic_vector(-6243,14),
		conv_std_logic_vector(-6239,14),
		conv_std_logic_vector(-6235,14),
		conv_std_logic_vector(-6231,14),
		conv_std_logic_vector(-6227,14),
		conv_std_logic_vector(-6223,14),
		conv_std_logic_vector(-6219,14),
		conv_std_logic_vector(-6215,14),
		conv_std_logic_vector(-6211,14),
		conv_std_logic_vector(-6207,14),
		conv_std_logic_vector(-6203,14),
		conv_std_logic_vector(-6198,14),
		conv_std_logic_vector(-6194,14),
		conv_std_logic_vector(-6190,14),
		conv_std_logic_vector(-6186,14),
		conv_std_logic_vector(-6182,14),
		conv_std_logic_vector(-6178,14),
		conv_std_logic_vector(-6174,14),
		conv_std_logic_vector(-6170,14),
		conv_std_logic_vector(-6165,14),
		conv_std_logic_vector(-6161,14),
		conv_std_logic_vector(-6157,14),
		conv_std_logic_vector(-6153,14),
		conv_std_logic_vector(-6149,14),
		conv_std_logic_vector(-6145,14),
		conv_std_logic_vector(-6141,14),
		conv_std_logic_vector(-6136,14),
		conv_std_logic_vector(-6132,14),
		conv_std_logic_vector(-6128,14),
		conv_std_logic_vector(-6124,14),
		conv_std_logic_vector(-6120,14),
		conv_std_logic_vector(-6116,14),
		conv_std_logic_vector(-6111,14),
		conv_std_logic_vector(-6107,14),
		conv_std_logic_vector(-6103,14),
		conv_std_logic_vector(-6099,14),
		conv_std_logic_vector(-6095,14),
		conv_std_logic_vector(-6090,14),
		conv_std_logic_vector(-6086,14),
		conv_std_logic_vector(-6082,14),
		conv_std_logic_vector(-6078,14),
		conv_std_logic_vector(-6074,14),
		conv_std_logic_vector(-6069,14),
		conv_std_logic_vector(-6065,14),
		conv_std_logic_vector(-6061,14),
		conv_std_logic_vector(-6057,14),
		conv_std_logic_vector(-6052,14),
		conv_std_logic_vector(-6048,14),
		conv_std_logic_vector(-6044,14),
		conv_std_logic_vector(-6040,14),
		conv_std_logic_vector(-6036,14),
		conv_std_logic_vector(-6031,14),
		conv_std_logic_vector(-6027,14),
		conv_std_logic_vector(-6023,14),
		conv_std_logic_vector(-6018,14),
		conv_std_logic_vector(-6014,14),
		conv_std_logic_vector(-6010,14),
		conv_std_logic_vector(-6006,14),
		conv_std_logic_vector(-6001,14),
		conv_std_logic_vector(-5997,14),
		conv_std_logic_vector(-5993,14),
		conv_std_logic_vector(-5989,14),
		conv_std_logic_vector(-5984,14),
		conv_std_logic_vector(-5980,14),
		conv_std_logic_vector(-5976,14),
		conv_std_logic_vector(-5971,14),
		conv_std_logic_vector(-5967,14),
		conv_std_logic_vector(-5963,14),
		conv_std_logic_vector(-5958,14),
		conv_std_logic_vector(-5954,14),
		conv_std_logic_vector(-5950,14),
		conv_std_logic_vector(-5946,14),
		conv_std_logic_vector(-5941,14),
		conv_std_logic_vector(-5937,14),
		conv_std_logic_vector(-5933,14),
		conv_std_logic_vector(-5928,14),
		conv_std_logic_vector(-5924,14),
		conv_std_logic_vector(-5920,14),
		conv_std_logic_vector(-5915,14),
		conv_std_logic_vector(-5911,14),
		conv_std_logic_vector(-5906,14),
		conv_std_logic_vector(-5902,14),
		conv_std_logic_vector(-5898,14),
		conv_std_logic_vector(-5893,14),
		conv_std_logic_vector(-5889,14),
		conv_std_logic_vector(-5885,14),
		conv_std_logic_vector(-5880,14),
		conv_std_logic_vector(-5876,14),
		conv_std_logic_vector(-5872,14),
		conv_std_logic_vector(-5867,14),
		conv_std_logic_vector(-5863,14),
		conv_std_logic_vector(-5858,14),
		conv_std_logic_vector(-5854,14),
		conv_std_logic_vector(-5850,14),
		conv_std_logic_vector(-5845,14),
		conv_std_logic_vector(-5841,14),
		conv_std_logic_vector(-5836,14),
		conv_std_logic_vector(-5832,14),
		conv_std_logic_vector(-5828,14),
		conv_std_logic_vector(-5823,14),
		conv_std_logic_vector(-5819,14),
		conv_std_logic_vector(-5814,14),
		conv_std_logic_vector(-5810,14),
		conv_std_logic_vector(-5805,14),
		conv_std_logic_vector(-5801,14),
		conv_std_logic_vector(-5797,14),
		conv_std_logic_vector(-5792,14),
		conv_std_logic_vector(-5788,14),
		conv_std_logic_vector(-5783,14),
		conv_std_logic_vector(-5779,14),
		conv_std_logic_vector(-5774,14),
		conv_std_logic_vector(-5770,14),
		conv_std_logic_vector(-5765,14),
		conv_std_logic_vector(-5761,14),
		conv_std_logic_vector(-5756,14),
		conv_std_logic_vector(-5752,14),
		conv_std_logic_vector(-5748,14),
		conv_std_logic_vector(-5743,14),
		conv_std_logic_vector(-5739,14),
		conv_std_logic_vector(-5734,14),
		conv_std_logic_vector(-5730,14),
		conv_std_logic_vector(-5725,14),
		conv_std_logic_vector(-5721,14),
		conv_std_logic_vector(-5716,14),
		conv_std_logic_vector(-5712,14),
		conv_std_logic_vector(-5707,14),
		conv_std_logic_vector(-5703,14),
		conv_std_logic_vector(-5698,14),
		conv_std_logic_vector(-5694,14),
		conv_std_logic_vector(-5689,14),
		conv_std_logic_vector(-5685,14),
		conv_std_logic_vector(-5680,14),
		conv_std_logic_vector(-5675,14),
		conv_std_logic_vector(-5671,14),
		conv_std_logic_vector(-5666,14),
		conv_std_logic_vector(-5662,14),
		conv_std_logic_vector(-5657,14),
		conv_std_logic_vector(-5653,14),
		conv_std_logic_vector(-5648,14),
		conv_std_logic_vector(-5644,14),
		conv_std_logic_vector(-5639,14),
		conv_std_logic_vector(-5635,14),
		conv_std_logic_vector(-5630,14),
		conv_std_logic_vector(-5625,14),
		conv_std_logic_vector(-5621,14),
		conv_std_logic_vector(-5616,14),
		conv_std_logic_vector(-5612,14),
		conv_std_logic_vector(-5607,14),
		conv_std_logic_vector(-5603,14),
		conv_std_logic_vector(-5598,14),
		conv_std_logic_vector(-5593,14),
		conv_std_logic_vector(-5589,14),
		conv_std_logic_vector(-5584,14),
		conv_std_logic_vector(-5580,14),
		conv_std_logic_vector(-5575,14),
		conv_std_logic_vector(-5570,14),
		conv_std_logic_vector(-5566,14),
		conv_std_logic_vector(-5561,14),
		conv_std_logic_vector(-5557,14),
		conv_std_logic_vector(-5552,14),
		conv_std_logic_vector(-5547,14),
		conv_std_logic_vector(-5543,14),
		conv_std_logic_vector(-5538,14),
		conv_std_logic_vector(-5533,14),
		conv_std_logic_vector(-5529,14),
		conv_std_logic_vector(-5524,14),
		conv_std_logic_vector(-5520,14),
		conv_std_logic_vector(-5515,14),
		conv_std_logic_vector(-5510,14),
		conv_std_logic_vector(-5506,14),
		conv_std_logic_vector(-5501,14),
		conv_std_logic_vector(-5496,14),
		conv_std_logic_vector(-5492,14),
		conv_std_logic_vector(-5487,14),
		conv_std_logic_vector(-5482,14),
		conv_std_logic_vector(-5478,14),
		conv_std_logic_vector(-5473,14),
		conv_std_logic_vector(-5468,14),
		conv_std_logic_vector(-5464,14),
		conv_std_logic_vector(-5459,14),
		conv_std_logic_vector(-5454,14),
		conv_std_logic_vector(-5450,14),
		conv_std_logic_vector(-5445,14),
		conv_std_logic_vector(-5440,14),
		conv_std_logic_vector(-5435,14),
		conv_std_logic_vector(-5431,14),
		conv_std_logic_vector(-5426,14),
		conv_std_logic_vector(-5421,14),
		conv_std_logic_vector(-5417,14),
		conv_std_logic_vector(-5412,14),
		conv_std_logic_vector(-5407,14),
		conv_std_logic_vector(-5402,14),
		conv_std_logic_vector(-5398,14),
		conv_std_logic_vector(-5393,14),
		conv_std_logic_vector(-5388,14),
		conv_std_logic_vector(-5384,14),
		conv_std_logic_vector(-5379,14),
		conv_std_logic_vector(-5374,14),
		conv_std_logic_vector(-5369,14),
		conv_std_logic_vector(-5365,14),
		conv_std_logic_vector(-5360,14),
		conv_std_logic_vector(-5355,14),
		conv_std_logic_vector(-5350,14),
		conv_std_logic_vector(-5346,14),
		conv_std_logic_vector(-5341,14),
		conv_std_logic_vector(-5336,14),
		conv_std_logic_vector(-5331,14),
		conv_std_logic_vector(-5326,14),
		conv_std_logic_vector(-5322,14),
		conv_std_logic_vector(-5317,14),
		conv_std_logic_vector(-5312,14),
		conv_std_logic_vector(-5307,14),
		conv_std_logic_vector(-5303,14),
		conv_std_logic_vector(-5298,14),
		conv_std_logic_vector(-5293,14),
		conv_std_logic_vector(-5288,14),
		conv_std_logic_vector(-5283,14),
		conv_std_logic_vector(-5279,14),
		conv_std_logic_vector(-5274,14),
		conv_std_logic_vector(-5269,14),
		conv_std_logic_vector(-5264,14),
		conv_std_logic_vector(-5259,14),
		conv_std_logic_vector(-5255,14),
		conv_std_logic_vector(-5250,14),
		conv_std_logic_vector(-5245,14),
		conv_std_logic_vector(-5240,14),
		conv_std_logic_vector(-5235,14),
		conv_std_logic_vector(-5230,14),
		conv_std_logic_vector(-5226,14),
		conv_std_logic_vector(-5221,14),
		conv_std_logic_vector(-5216,14),
		conv_std_logic_vector(-5211,14),
		conv_std_logic_vector(-5206,14),
		conv_std_logic_vector(-5201,14),
		conv_std_logic_vector(-5196,14),
		conv_std_logic_vector(-5192,14),
		conv_std_logic_vector(-5187,14),
		conv_std_logic_vector(-5182,14),
		conv_std_logic_vector(-5177,14),
		conv_std_logic_vector(-5172,14),
		conv_std_logic_vector(-5167,14),
		conv_std_logic_vector(-5162,14),
		conv_std_logic_vector(-5157,14),
		conv_std_logic_vector(-5153,14),
		conv_std_logic_vector(-5148,14),
		conv_std_logic_vector(-5143,14),
		conv_std_logic_vector(-5138,14),
		conv_std_logic_vector(-5133,14),
		conv_std_logic_vector(-5128,14),
		conv_std_logic_vector(-5123,14),
		conv_std_logic_vector(-5118,14),
		conv_std_logic_vector(-5113,14),
		conv_std_logic_vector(-5109,14),
		conv_std_logic_vector(-5104,14),
		conv_std_logic_vector(-5099,14),
		conv_std_logic_vector(-5094,14),
		conv_std_logic_vector(-5089,14),
		conv_std_logic_vector(-5084,14),
		conv_std_logic_vector(-5079,14),
		conv_std_logic_vector(-5074,14),
		conv_std_logic_vector(-5069,14),
		conv_std_logic_vector(-5064,14),
		conv_std_logic_vector(-5059,14),
		conv_std_logic_vector(-5054,14),
		conv_std_logic_vector(-5049,14),
		conv_std_logic_vector(-5044,14),
		conv_std_logic_vector(-5039,14),
		conv_std_logic_vector(-5035,14),
		conv_std_logic_vector(-5030,14),
		conv_std_logic_vector(-5025,14),
		conv_std_logic_vector(-5020,14),
		conv_std_logic_vector(-5015,14),
		conv_std_logic_vector(-5010,14),
		conv_std_logic_vector(-5005,14),
		conv_std_logic_vector(-5000,14),
		conv_std_logic_vector(-4995,14),
		conv_std_logic_vector(-4990,14),
		conv_std_logic_vector(-4985,14),
		conv_std_logic_vector(-4980,14),
		conv_std_logic_vector(-4975,14),
		conv_std_logic_vector(-4970,14),
		conv_std_logic_vector(-4965,14),
		conv_std_logic_vector(-4960,14),
		conv_std_logic_vector(-4955,14),
		conv_std_logic_vector(-4950,14),
		conv_std_logic_vector(-4945,14),
		conv_std_logic_vector(-4940,14),
		conv_std_logic_vector(-4935,14),
		conv_std_logic_vector(-4930,14),
		conv_std_logic_vector(-4925,14),
		conv_std_logic_vector(-4920,14),
		conv_std_logic_vector(-4915,14),
		conv_std_logic_vector(-4910,14),
		conv_std_logic_vector(-4905,14),
		conv_std_logic_vector(-4900,14),
		conv_std_logic_vector(-4895,14),
		conv_std_logic_vector(-4890,14),
		conv_std_logic_vector(-4885,14),
		conv_std_logic_vector(-4879,14),
		conv_std_logic_vector(-4874,14),
		conv_std_logic_vector(-4869,14),
		conv_std_logic_vector(-4864,14),
		conv_std_logic_vector(-4859,14),
		conv_std_logic_vector(-4854,14),
		conv_std_logic_vector(-4849,14),
		conv_std_logic_vector(-4844,14),
		conv_std_logic_vector(-4839,14),
		conv_std_logic_vector(-4834,14),
		conv_std_logic_vector(-4829,14),
		conv_std_logic_vector(-4824,14),
		conv_std_logic_vector(-4819,14),
		conv_std_logic_vector(-4814,14),
		conv_std_logic_vector(-4809,14),
		conv_std_logic_vector(-4803,14),
		conv_std_logic_vector(-4798,14),
		conv_std_logic_vector(-4793,14),
		conv_std_logic_vector(-4788,14),
		conv_std_logic_vector(-4783,14),
		conv_std_logic_vector(-4778,14),
		conv_std_logic_vector(-4773,14),
		conv_std_logic_vector(-4768,14),
		conv_std_logic_vector(-4763,14),
		conv_std_logic_vector(-4758,14),
		conv_std_logic_vector(-4752,14),
		conv_std_logic_vector(-4747,14),
		conv_std_logic_vector(-4742,14),
		conv_std_logic_vector(-4737,14),
		conv_std_logic_vector(-4732,14),
		conv_std_logic_vector(-4727,14),
		conv_std_logic_vector(-4722,14),
		conv_std_logic_vector(-4717,14),
		conv_std_logic_vector(-4711,14),
		conv_std_logic_vector(-4706,14),
		conv_std_logic_vector(-4701,14),
		conv_std_logic_vector(-4696,14),
		conv_std_logic_vector(-4691,14),
		conv_std_logic_vector(-4686,14),
		conv_std_logic_vector(-4680,14),
		conv_std_logic_vector(-4675,14),
		conv_std_logic_vector(-4670,14),
		conv_std_logic_vector(-4665,14),
		conv_std_logic_vector(-4660,14),
		conv_std_logic_vector(-4655,14),
		conv_std_logic_vector(-4650,14),
		conv_std_logic_vector(-4644,14),
		conv_std_logic_vector(-4639,14),
		conv_std_logic_vector(-4634,14),
		conv_std_logic_vector(-4629,14),
		conv_std_logic_vector(-4624,14),
		conv_std_logic_vector(-4618,14),
		conv_std_logic_vector(-4613,14),
		conv_std_logic_vector(-4608,14),
		conv_std_logic_vector(-4603,14),
		conv_std_logic_vector(-4598,14),
		conv_std_logic_vector(-4592,14),
		conv_std_logic_vector(-4587,14),
		conv_std_logic_vector(-4582,14),
		conv_std_logic_vector(-4577,14),
		conv_std_logic_vector(-4572,14),
		conv_std_logic_vector(-4566,14),
		conv_std_logic_vector(-4561,14),
		conv_std_logic_vector(-4556,14),
		conv_std_logic_vector(-4551,14),
		conv_std_logic_vector(-4546,14),
		conv_std_logic_vector(-4540,14),
		conv_std_logic_vector(-4535,14),
		conv_std_logic_vector(-4530,14),
		conv_std_logic_vector(-4525,14),
		conv_std_logic_vector(-4519,14),
		conv_std_logic_vector(-4514,14),
		conv_std_logic_vector(-4509,14),
		conv_std_logic_vector(-4504,14),
		conv_std_logic_vector(-4498,14),
		conv_std_logic_vector(-4493,14),
		conv_std_logic_vector(-4488,14),
		conv_std_logic_vector(-4483,14),
		conv_std_logic_vector(-4477,14),
		conv_std_logic_vector(-4472,14),
		conv_std_logic_vector(-4467,14),
		conv_std_logic_vector(-4462,14),
		conv_std_logic_vector(-4456,14),
		conv_std_logic_vector(-4451,14),
		conv_std_logic_vector(-4446,14),
		conv_std_logic_vector(-4440,14),
		conv_std_logic_vector(-4435,14),
		conv_std_logic_vector(-4430,14),
		conv_std_logic_vector(-4425,14),
		conv_std_logic_vector(-4419,14),
		conv_std_logic_vector(-4414,14),
		conv_std_logic_vector(-4409,14),
		conv_std_logic_vector(-4403,14),
		conv_std_logic_vector(-4398,14),
		conv_std_logic_vector(-4393,14),
		conv_std_logic_vector(-4388,14),
		conv_std_logic_vector(-4382,14),
		conv_std_logic_vector(-4377,14),
		conv_std_logic_vector(-4372,14),
		conv_std_logic_vector(-4366,14),
		conv_std_logic_vector(-4361,14),
		conv_std_logic_vector(-4356,14),
		conv_std_logic_vector(-4350,14),
		conv_std_logic_vector(-4345,14),
		conv_std_logic_vector(-4340,14),
		conv_std_logic_vector(-4334,14),
		conv_std_logic_vector(-4329,14),
		conv_std_logic_vector(-4324,14),
		conv_std_logic_vector(-4318,14),
		conv_std_logic_vector(-4313,14),
		conv_std_logic_vector(-4308,14),
		conv_std_logic_vector(-4302,14),
		conv_std_logic_vector(-4297,14),
		conv_std_logic_vector(-4292,14),
		conv_std_logic_vector(-4286,14),
		conv_std_logic_vector(-4281,14),
		conv_std_logic_vector(-4276,14),
		conv_std_logic_vector(-4270,14),
		conv_std_logic_vector(-4265,14),
		conv_std_logic_vector(-4259,14),
		conv_std_logic_vector(-4254,14),
		conv_std_logic_vector(-4249,14),
		conv_std_logic_vector(-4243,14),
		conv_std_logic_vector(-4238,14),
		conv_std_logic_vector(-4233,14),
		conv_std_logic_vector(-4227,14),
		conv_std_logic_vector(-4222,14),
		conv_std_logic_vector(-4216,14),
		conv_std_logic_vector(-4211,14),
		conv_std_logic_vector(-4206,14),
		conv_std_logic_vector(-4200,14),
		conv_std_logic_vector(-4195,14),
		conv_std_logic_vector(-4189,14),
		conv_std_logic_vector(-4184,14),
		conv_std_logic_vector(-4179,14),
		conv_std_logic_vector(-4173,14),
		conv_std_logic_vector(-4168,14),
		conv_std_logic_vector(-4162,14),
		conv_std_logic_vector(-4157,14),
		conv_std_logic_vector(-4152,14),
		conv_std_logic_vector(-4146,14),
		conv_std_logic_vector(-4141,14),
		conv_std_logic_vector(-4135,14),
		conv_std_logic_vector(-4130,14),
		conv_std_logic_vector(-4124,14),
		conv_std_logic_vector(-4119,14),
		conv_std_logic_vector(-4114,14),
		conv_std_logic_vector(-4108,14),
		conv_std_logic_vector(-4103,14),
		conv_std_logic_vector(-4097,14),
		conv_std_logic_vector(-4092,14),
		conv_std_logic_vector(-4086,14),
		conv_std_logic_vector(-4081,14),
		conv_std_logic_vector(-4076,14),
		conv_std_logic_vector(-4070,14),
		conv_std_logic_vector(-4065,14),
		conv_std_logic_vector(-4059,14),
		conv_std_logic_vector(-4054,14),
		conv_std_logic_vector(-4048,14),
		conv_std_logic_vector(-4043,14),
		conv_std_logic_vector(-4037,14),
		conv_std_logic_vector(-4032,14),
		conv_std_logic_vector(-4026,14),
		conv_std_logic_vector(-4021,14),
		conv_std_logic_vector(-4015,14),
		conv_std_logic_vector(-4010,14),
		conv_std_logic_vector(-4004,14),
		conv_std_logic_vector(-3999,14),
		conv_std_logic_vector(-3994,14),
		conv_std_logic_vector(-3988,14),
		conv_std_logic_vector(-3983,14),
		conv_std_logic_vector(-3977,14),
		conv_std_logic_vector(-3972,14),
		conv_std_logic_vector(-3966,14),
		conv_std_logic_vector(-3961,14),
		conv_std_logic_vector(-3955,14),
		conv_std_logic_vector(-3950,14),
		conv_std_logic_vector(-3944,14),
		conv_std_logic_vector(-3939,14),
		conv_std_logic_vector(-3933,14),
		conv_std_logic_vector(-3928,14),
		conv_std_logic_vector(-3922,14),
		conv_std_logic_vector(-3916,14),
		conv_std_logic_vector(-3911,14),
		conv_std_logic_vector(-3905,14),
		conv_std_logic_vector(-3900,14),
		conv_std_logic_vector(-3894,14),
		conv_std_logic_vector(-3889,14),
		conv_std_logic_vector(-3883,14),
		conv_std_logic_vector(-3878,14),
		conv_std_logic_vector(-3872,14),
		conv_std_logic_vector(-3867,14),
		conv_std_logic_vector(-3861,14),
		conv_std_logic_vector(-3856,14),
		conv_std_logic_vector(-3850,14),
		conv_std_logic_vector(-3845,14),
		conv_std_logic_vector(-3839,14),
		conv_std_logic_vector(-3833,14),
		conv_std_logic_vector(-3828,14),
		conv_std_logic_vector(-3822,14),
		conv_std_logic_vector(-3817,14),
		conv_std_logic_vector(-3811,14),
		conv_std_logic_vector(-3806,14),
		conv_std_logic_vector(-3800,14),
		conv_std_logic_vector(-3795,14),
		conv_std_logic_vector(-3789,14),
		conv_std_logic_vector(-3783,14),
		conv_std_logic_vector(-3778,14),
		conv_std_logic_vector(-3772,14),
		conv_std_logic_vector(-3767,14),
		conv_std_logic_vector(-3761,14),
		conv_std_logic_vector(-3755,14),
		conv_std_logic_vector(-3750,14),
		conv_std_logic_vector(-3744,14),
		conv_std_logic_vector(-3739,14),
		conv_std_logic_vector(-3733,14),
		conv_std_logic_vector(-3728,14),
		conv_std_logic_vector(-3722,14),
		conv_std_logic_vector(-3716,14),
		conv_std_logic_vector(-3711,14),
		conv_std_logic_vector(-3705,14),
		conv_std_logic_vector(-3700,14),
		conv_std_logic_vector(-3694,14),
		conv_std_logic_vector(-3688,14),
		conv_std_logic_vector(-3683,14),
		conv_std_logic_vector(-3677,14),
		conv_std_logic_vector(-3671,14),
		conv_std_logic_vector(-3666,14),
		conv_std_logic_vector(-3660,14),
		conv_std_logic_vector(-3655,14),
		conv_std_logic_vector(-3649,14),
		conv_std_logic_vector(-3643,14),
		conv_std_logic_vector(-3638,14),
		conv_std_logic_vector(-3632,14),
		conv_std_logic_vector(-3626,14),
		conv_std_logic_vector(-3621,14),
		conv_std_logic_vector(-3615,14),
		conv_std_logic_vector(-3610,14),
		conv_std_logic_vector(-3604,14),
		conv_std_logic_vector(-3598,14),
		conv_std_logic_vector(-3593,14),
		conv_std_logic_vector(-3587,14),
		conv_std_logic_vector(-3581,14),
		conv_std_logic_vector(-3576,14),
		conv_std_logic_vector(-3570,14),
		conv_std_logic_vector(-3564,14),
		conv_std_logic_vector(-3559,14),
		conv_std_logic_vector(-3553,14),
		conv_std_logic_vector(-3547,14),
		conv_std_logic_vector(-3542,14),
		conv_std_logic_vector(-3536,14),
		conv_std_logic_vector(-3530,14),
		conv_std_logic_vector(-3525,14),
		conv_std_logic_vector(-3519,14),
		conv_std_logic_vector(-3513,14),
		conv_std_logic_vector(-3508,14),
		conv_std_logic_vector(-3502,14),
		conv_std_logic_vector(-3496,14),
		conv_std_logic_vector(-3491,14),
		conv_std_logic_vector(-3485,14),
		conv_std_logic_vector(-3479,14),
		conv_std_logic_vector(-3474,14),
		conv_std_logic_vector(-3468,14),
		conv_std_logic_vector(-3462,14),
		conv_std_logic_vector(-3457,14),
		conv_std_logic_vector(-3451,14),
		conv_std_logic_vector(-3445,14),
		conv_std_logic_vector(-3439,14),
		conv_std_logic_vector(-3434,14),
		conv_std_logic_vector(-3428,14),
		conv_std_logic_vector(-3422,14),
		conv_std_logic_vector(-3417,14),
		conv_std_logic_vector(-3411,14),
		conv_std_logic_vector(-3405,14),
		conv_std_logic_vector(-3399,14),
		conv_std_logic_vector(-3394,14),
		conv_std_logic_vector(-3388,14),
		conv_std_logic_vector(-3382,14),
		conv_std_logic_vector(-3377,14),
		conv_std_logic_vector(-3371,14),
		conv_std_logic_vector(-3365,14),
		conv_std_logic_vector(-3359,14),
		conv_std_logic_vector(-3354,14),
		conv_std_logic_vector(-3348,14),
		conv_std_logic_vector(-3342,14),
		conv_std_logic_vector(-3336,14),
		conv_std_logic_vector(-3331,14),
		conv_std_logic_vector(-3325,14),
		conv_std_logic_vector(-3319,14),
		conv_std_logic_vector(-3313,14),
		conv_std_logic_vector(-3308,14),
		conv_std_logic_vector(-3302,14),
		conv_std_logic_vector(-3296,14),
		conv_std_logic_vector(-3290,14),
		conv_std_logic_vector(-3285,14),
		conv_std_logic_vector(-3279,14),
		conv_std_logic_vector(-3273,14),
		conv_std_logic_vector(-3267,14),
		conv_std_logic_vector(-3262,14),
		conv_std_logic_vector(-3256,14),
		conv_std_logic_vector(-3250,14),
		conv_std_logic_vector(-3244,14),
		conv_std_logic_vector(-3239,14),
		conv_std_logic_vector(-3233,14),
		conv_std_logic_vector(-3227,14),
		conv_std_logic_vector(-3221,14),
		conv_std_logic_vector(-3216,14),
		conv_std_logic_vector(-3210,14),
		conv_std_logic_vector(-3204,14),
		conv_std_logic_vector(-3198,14),
		conv_std_logic_vector(-3192,14),
		conv_std_logic_vector(-3187,14),
		conv_std_logic_vector(-3181,14),
		conv_std_logic_vector(-3175,14),
		conv_std_logic_vector(-3169,14),
		conv_std_logic_vector(-3163,14),
		conv_std_logic_vector(-3158,14),
		conv_std_logic_vector(-3152,14),
		conv_std_logic_vector(-3146,14),
		conv_std_logic_vector(-3140,14),
		conv_std_logic_vector(-3134,14),
		conv_std_logic_vector(-3129,14),
		conv_std_logic_vector(-3123,14),
		conv_std_logic_vector(-3117,14),
		conv_std_logic_vector(-3111,14),
		conv_std_logic_vector(-3105,14),
		conv_std_logic_vector(-3100,14),
		conv_std_logic_vector(-3094,14),
		conv_std_logic_vector(-3088,14),
		conv_std_logic_vector(-3082,14),
		conv_std_logic_vector(-3076,14),
		conv_std_logic_vector(-3070,14),
		conv_std_logic_vector(-3065,14),
		conv_std_logic_vector(-3059,14),
		conv_std_logic_vector(-3053,14),
		conv_std_logic_vector(-3047,14),
		conv_std_logic_vector(-3041,14),
		conv_std_logic_vector(-3035,14),
		conv_std_logic_vector(-3030,14),
		conv_std_logic_vector(-3024,14),
		conv_std_logic_vector(-3018,14),
		conv_std_logic_vector(-3012,14),
		conv_std_logic_vector(-3006,14),
		conv_std_logic_vector(-3000,14),
		conv_std_logic_vector(-2995,14),
		conv_std_logic_vector(-2989,14),
		conv_std_logic_vector(-2983,14),
		conv_std_logic_vector(-2977,14),
		conv_std_logic_vector(-2971,14),
		conv_std_logic_vector(-2965,14),
		conv_std_logic_vector(-2959,14),
		conv_std_logic_vector(-2954,14),
		conv_std_logic_vector(-2948,14),
		conv_std_logic_vector(-2942,14),
		conv_std_logic_vector(-2936,14),
		conv_std_logic_vector(-2930,14),
		conv_std_logic_vector(-2924,14),
		conv_std_logic_vector(-2918,14),
		conv_std_logic_vector(-2913,14),
		conv_std_logic_vector(-2907,14),
		conv_std_logic_vector(-2901,14),
		conv_std_logic_vector(-2895,14),
		conv_std_logic_vector(-2889,14),
		conv_std_logic_vector(-2883,14),
		conv_std_logic_vector(-2877,14),
		conv_std_logic_vector(-2871,14),
		conv_std_logic_vector(-2866,14),
		conv_std_logic_vector(-2860,14),
		conv_std_logic_vector(-2854,14),
		conv_std_logic_vector(-2848,14),
		conv_std_logic_vector(-2842,14),
		conv_std_logic_vector(-2836,14),
		conv_std_logic_vector(-2830,14),
		conv_std_logic_vector(-2824,14),
		conv_std_logic_vector(-2818,14),
		conv_std_logic_vector(-2812,14),
		conv_std_logic_vector(-2807,14),
		conv_std_logic_vector(-2801,14),
		conv_std_logic_vector(-2795,14),
		conv_std_logic_vector(-2789,14),
		conv_std_logic_vector(-2783,14),
		conv_std_logic_vector(-2777,14),
		conv_std_logic_vector(-2771,14),
		conv_std_logic_vector(-2765,14),
		conv_std_logic_vector(-2759,14),
		conv_std_logic_vector(-2753,14),
		conv_std_logic_vector(-2747,14),
		conv_std_logic_vector(-2742,14),
		conv_std_logic_vector(-2736,14),
		conv_std_logic_vector(-2730,14),
		conv_std_logic_vector(-2724,14),
		conv_std_logic_vector(-2718,14),
		conv_std_logic_vector(-2712,14),
		conv_std_logic_vector(-2706,14),
		conv_std_logic_vector(-2700,14),
		conv_std_logic_vector(-2694,14),
		conv_std_logic_vector(-2688,14),
		conv_std_logic_vector(-2682,14),
		conv_std_logic_vector(-2676,14),
		conv_std_logic_vector(-2670,14),
		conv_std_logic_vector(-2664,14),
		conv_std_logic_vector(-2658,14),
		conv_std_logic_vector(-2653,14),
		conv_std_logic_vector(-2647,14),
		conv_std_logic_vector(-2641,14),
		conv_std_logic_vector(-2635,14),
		conv_std_logic_vector(-2629,14),
		conv_std_logic_vector(-2623,14),
		conv_std_logic_vector(-2617,14),
		conv_std_logic_vector(-2611,14),
		conv_std_logic_vector(-2605,14),
		conv_std_logic_vector(-2599,14),
		conv_std_logic_vector(-2593,14),
		conv_std_logic_vector(-2587,14),
		conv_std_logic_vector(-2581,14),
		conv_std_logic_vector(-2575,14),
		conv_std_logic_vector(-2569,14),
		conv_std_logic_vector(-2563,14),
		conv_std_logic_vector(-2557,14),
		conv_std_logic_vector(-2551,14),
		conv_std_logic_vector(-2545,14),
		conv_std_logic_vector(-2539,14),
		conv_std_logic_vector(-2533,14),
		conv_std_logic_vector(-2527,14),
		conv_std_logic_vector(-2521,14),
		conv_std_logic_vector(-2515,14),
		conv_std_logic_vector(-2509,14),
		conv_std_logic_vector(-2503,14),
		conv_std_logic_vector(-2497,14),
		conv_std_logic_vector(-2491,14),
		conv_std_logic_vector(-2486,14),
		conv_std_logic_vector(-2480,14),
		conv_std_logic_vector(-2474,14),
		conv_std_logic_vector(-2468,14),
		conv_std_logic_vector(-2462,14),
		conv_std_logic_vector(-2456,14),
		conv_std_logic_vector(-2450,14),
		conv_std_logic_vector(-2444,14),
		conv_std_logic_vector(-2438,14),
		conv_std_logic_vector(-2432,14),
		conv_std_logic_vector(-2426,14),
		conv_std_logic_vector(-2420,14),
		conv_std_logic_vector(-2414,14),
		conv_std_logic_vector(-2408,14),
		conv_std_logic_vector(-2402,14),
		conv_std_logic_vector(-2396,14),
		conv_std_logic_vector(-2390,14),
		conv_std_logic_vector(-2384,14),
		conv_std_logic_vector(-2378,14),
		conv_std_logic_vector(-2371,14),
		conv_std_logic_vector(-2365,14),
		conv_std_logic_vector(-2359,14),
		conv_std_logic_vector(-2353,14),
		conv_std_logic_vector(-2347,14),
		conv_std_logic_vector(-2341,14),
		conv_std_logic_vector(-2335,14),
		conv_std_logic_vector(-2329,14),
		conv_std_logic_vector(-2323,14),
		conv_std_logic_vector(-2317,14),
		conv_std_logic_vector(-2311,14),
		conv_std_logic_vector(-2305,14),
		conv_std_logic_vector(-2299,14),
		conv_std_logic_vector(-2293,14),
		conv_std_logic_vector(-2287,14),
		conv_std_logic_vector(-2281,14),
		conv_std_logic_vector(-2275,14),
		conv_std_logic_vector(-2269,14),
		conv_std_logic_vector(-2263,14),
		conv_std_logic_vector(-2257,14),
		conv_std_logic_vector(-2251,14),
		conv_std_logic_vector(-2245,14),
		conv_std_logic_vector(-2239,14),
		conv_std_logic_vector(-2233,14),
		conv_std_logic_vector(-2227,14),
		conv_std_logic_vector(-2221,14),
		conv_std_logic_vector(-2215,14),
		conv_std_logic_vector(-2209,14),
		conv_std_logic_vector(-2203,14),
		conv_std_logic_vector(-2197,14),
		conv_std_logic_vector(-2190,14),
		conv_std_logic_vector(-2184,14),
		conv_std_logic_vector(-2178,14),
		conv_std_logic_vector(-2172,14),
		conv_std_logic_vector(-2166,14),
		conv_std_logic_vector(-2160,14),
		conv_std_logic_vector(-2154,14),
		conv_std_logic_vector(-2148,14),
		conv_std_logic_vector(-2142,14),
		conv_std_logic_vector(-2136,14),
		conv_std_logic_vector(-2130,14),
		conv_std_logic_vector(-2124,14),
		conv_std_logic_vector(-2118,14),
		conv_std_logic_vector(-2112,14),
		conv_std_logic_vector(-2106,14),
		conv_std_logic_vector(-2100,14),
		conv_std_logic_vector(-2093,14),
		conv_std_logic_vector(-2087,14),
		conv_std_logic_vector(-2081,14),
		conv_std_logic_vector(-2075,14),
		conv_std_logic_vector(-2069,14),
		conv_std_logic_vector(-2063,14),
		conv_std_logic_vector(-2057,14),
		conv_std_logic_vector(-2051,14),
		conv_std_logic_vector(-2045,14),
		conv_std_logic_vector(-2039,14),
		conv_std_logic_vector(-2033,14),
		conv_std_logic_vector(-2027,14),
		conv_std_logic_vector(-2020,14),
		conv_std_logic_vector(-2014,14),
		conv_std_logic_vector(-2008,14),
		conv_std_logic_vector(-2002,14),
		conv_std_logic_vector(-1996,14),
		conv_std_logic_vector(-1990,14),
		conv_std_logic_vector(-1984,14),
		conv_std_logic_vector(-1978,14),
		conv_std_logic_vector(-1972,14),
		conv_std_logic_vector(-1966,14),
		conv_std_logic_vector(-1960,14),
		conv_std_logic_vector(-1953,14),
		conv_std_logic_vector(-1947,14),
		conv_std_logic_vector(-1941,14),
		conv_std_logic_vector(-1935,14),
		conv_std_logic_vector(-1929,14),
		conv_std_logic_vector(-1923,14),
		conv_std_logic_vector(-1917,14),
		conv_std_logic_vector(-1911,14),
		conv_std_logic_vector(-1905,14),
		conv_std_logic_vector(-1898,14),
		conv_std_logic_vector(-1892,14),
		conv_std_logic_vector(-1886,14),
		conv_std_logic_vector(-1880,14),
		conv_std_logic_vector(-1874,14),
		conv_std_logic_vector(-1868,14),
		conv_std_logic_vector(-1862,14),
		conv_std_logic_vector(-1856,14),
		conv_std_logic_vector(-1850,14),
		conv_std_logic_vector(-1843,14),
		conv_std_logic_vector(-1837,14),
		conv_std_logic_vector(-1831,14),
		conv_std_logic_vector(-1825,14),
		conv_std_logic_vector(-1819,14),
		conv_std_logic_vector(-1813,14),
		conv_std_logic_vector(-1807,14),
		conv_std_logic_vector(-1801,14),
		conv_std_logic_vector(-1794,14),
		conv_std_logic_vector(-1788,14),
		conv_std_logic_vector(-1782,14),
		conv_std_logic_vector(-1776,14),
		conv_std_logic_vector(-1770,14),
		conv_std_logic_vector(-1764,14),
		conv_std_logic_vector(-1758,14),
		conv_std_logic_vector(-1751,14),
		conv_std_logic_vector(-1745,14),
		conv_std_logic_vector(-1739,14),
		conv_std_logic_vector(-1733,14),
		conv_std_logic_vector(-1727,14),
		conv_std_logic_vector(-1721,14),
		conv_std_logic_vector(-1715,14),
		conv_std_logic_vector(-1708,14),
		conv_std_logic_vector(-1702,14),
		conv_std_logic_vector(-1696,14),
		conv_std_logic_vector(-1690,14),
		conv_std_logic_vector(-1684,14),
		conv_std_logic_vector(-1678,14),
		conv_std_logic_vector(-1672,14),
		conv_std_logic_vector(-1665,14),
		conv_std_logic_vector(-1659,14),
		conv_std_logic_vector(-1653,14),
		conv_std_logic_vector(-1647,14),
		conv_std_logic_vector(-1641,14),
		conv_std_logic_vector(-1635,14),
		conv_std_logic_vector(-1628,14),
		conv_std_logic_vector(-1622,14),
		conv_std_logic_vector(-1616,14),
		conv_std_logic_vector(-1610,14),
		conv_std_logic_vector(-1604,14),
		conv_std_logic_vector(-1598,14),
		conv_std_logic_vector(-1592,14),
		conv_std_logic_vector(-1585,14),
		conv_std_logic_vector(-1579,14),
		conv_std_logic_vector(-1573,14),
		conv_std_logic_vector(-1567,14),
		conv_std_logic_vector(-1561,14),
		conv_std_logic_vector(-1555,14),
		conv_std_logic_vector(-1548,14),
		conv_std_logic_vector(-1542,14),
		conv_std_logic_vector(-1536,14),
		conv_std_logic_vector(-1530,14),
		conv_std_logic_vector(-1524,14),
		conv_std_logic_vector(-1517,14),
		conv_std_logic_vector(-1511,14),
		conv_std_logic_vector(-1505,14),
		conv_std_logic_vector(-1499,14),
		conv_std_logic_vector(-1493,14),
		conv_std_logic_vector(-1487,14),
		conv_std_logic_vector(-1480,14),
		conv_std_logic_vector(-1474,14),
		conv_std_logic_vector(-1468,14),
		conv_std_logic_vector(-1462,14),
		conv_std_logic_vector(-1456,14),
		conv_std_logic_vector(-1450,14),
		conv_std_logic_vector(-1443,14),
		conv_std_logic_vector(-1437,14),
		conv_std_logic_vector(-1431,14),
		conv_std_logic_vector(-1425,14),
		conv_std_logic_vector(-1419,14),
		conv_std_logic_vector(-1412,14),
		conv_std_logic_vector(-1406,14),
		conv_std_logic_vector(-1400,14),
		conv_std_logic_vector(-1394,14),
		conv_std_logic_vector(-1388,14),
		conv_std_logic_vector(-1381,14),
		conv_std_logic_vector(-1375,14),
		conv_std_logic_vector(-1369,14),
		conv_std_logic_vector(-1363,14),
		conv_std_logic_vector(-1357,14),
		conv_std_logic_vector(-1350,14),
		conv_std_logic_vector(-1344,14),
		conv_std_logic_vector(-1338,14),
		conv_std_logic_vector(-1332,14),
		conv_std_logic_vector(-1326,14),
		conv_std_logic_vector(-1319,14),
		conv_std_logic_vector(-1313,14),
		conv_std_logic_vector(-1307,14),
		conv_std_logic_vector(-1301,14),
		conv_std_logic_vector(-1295,14),
		conv_std_logic_vector(-1288,14),
		conv_std_logic_vector(-1282,14),
		conv_std_logic_vector(-1276,14),
		conv_std_logic_vector(-1270,14),
		conv_std_logic_vector(-1264,14),
		conv_std_logic_vector(-1257,14),
		conv_std_logic_vector(-1251,14),
		conv_std_logic_vector(-1245,14),
		conv_std_logic_vector(-1239,14),
		conv_std_logic_vector(-1233,14),
		conv_std_logic_vector(-1226,14),
		conv_std_logic_vector(-1220,14),
		conv_std_logic_vector(-1214,14),
		conv_std_logic_vector(-1208,14),
		conv_std_logic_vector(-1202,14),
		conv_std_logic_vector(-1195,14),
		conv_std_logic_vector(-1189,14),
		conv_std_logic_vector(-1183,14),
		conv_std_logic_vector(-1177,14),
		conv_std_logic_vector(-1170,14),
		conv_std_logic_vector(-1164,14),
		conv_std_logic_vector(-1158,14),
		conv_std_logic_vector(-1152,14),
		conv_std_logic_vector(-1146,14),
		conv_std_logic_vector(-1139,14),
		conv_std_logic_vector(-1133,14),
		conv_std_logic_vector(-1127,14),
		conv_std_logic_vector(-1121,14),
		conv_std_logic_vector(-1114,14),
		conv_std_logic_vector(-1108,14),
		conv_std_logic_vector(-1102,14),
		conv_std_logic_vector(-1096,14),
		conv_std_logic_vector(-1090,14),
		conv_std_logic_vector(-1083,14),
		conv_std_logic_vector(-1077,14),
		conv_std_logic_vector(-1071,14),
		conv_std_logic_vector(-1065,14),
		conv_std_logic_vector(-1058,14),
		conv_std_logic_vector(-1052,14),
		conv_std_logic_vector(-1046,14),
		conv_std_logic_vector(-1040,14),
		conv_std_logic_vector(-1033,14),
		conv_std_logic_vector(-1027,14),
		conv_std_logic_vector(-1021,14),
		conv_std_logic_vector(-1015,14),
		conv_std_logic_vector(-1009,14),
		conv_std_logic_vector(-1002,14),
		conv_std_logic_vector(-996,14),
		conv_std_logic_vector(-990,14),
		conv_std_logic_vector(-984,14),
		conv_std_logic_vector(-977,14),
		conv_std_logic_vector(-971,14),
		conv_std_logic_vector(-965,14),
		conv_std_logic_vector(-959,14),
		conv_std_logic_vector(-952,14),
		conv_std_logic_vector(-946,14),
		conv_std_logic_vector(-940,14),
		conv_std_logic_vector(-934,14),
		conv_std_logic_vector(-927,14),
		conv_std_logic_vector(-921,14),
		conv_std_logic_vector(-915,14),
		conv_std_logic_vector(-909,14),
		conv_std_logic_vector(-902,14),
		conv_std_logic_vector(-896,14),
		conv_std_logic_vector(-890,14),
		conv_std_logic_vector(-884,14),
		conv_std_logic_vector(-877,14),
		conv_std_logic_vector(-871,14),
		conv_std_logic_vector(-865,14),
		conv_std_logic_vector(-859,14),
		conv_std_logic_vector(-852,14),
		conv_std_logic_vector(-846,14),
		conv_std_logic_vector(-840,14),
		conv_std_logic_vector(-834,14),
		conv_std_logic_vector(-827,14),
		conv_std_logic_vector(-821,14),
		conv_std_logic_vector(-815,14),
		conv_std_logic_vector(-809,14),
		conv_std_logic_vector(-802,14),
		conv_std_logic_vector(-796,14),
		conv_std_logic_vector(-790,14),
		conv_std_logic_vector(-784,14),
		conv_std_logic_vector(-777,14),
		conv_std_logic_vector(-771,14),
		conv_std_logic_vector(-765,14),
		conv_std_logic_vector(-759,14),
		conv_std_logic_vector(-752,14),
		conv_std_logic_vector(-746,14),
		conv_std_logic_vector(-740,14),
		conv_std_logic_vector(-734,14),
		conv_std_logic_vector(-727,14),
		conv_std_logic_vector(-721,14),
		conv_std_logic_vector(-715,14),
		conv_std_logic_vector(-709,14),
		conv_std_logic_vector(-702,14),
		conv_std_logic_vector(-696,14),
		conv_std_logic_vector(-690,14),
		conv_std_logic_vector(-684,14),
		conv_std_logic_vector(-677,14),
		conv_std_logic_vector(-671,14),
		conv_std_logic_vector(-665,14),
		conv_std_logic_vector(-659,14),
		conv_std_logic_vector(-652,14),
		conv_std_logic_vector(-646,14),
		conv_std_logic_vector(-640,14),
		conv_std_logic_vector(-633,14),
		conv_std_logic_vector(-627,14),
		conv_std_logic_vector(-621,14),
		conv_std_logic_vector(-615,14),
		conv_std_logic_vector(-608,14),
		conv_std_logic_vector(-602,14),
		conv_std_logic_vector(-596,14),
		conv_std_logic_vector(-590,14),
		conv_std_logic_vector(-583,14),
		conv_std_logic_vector(-577,14),
		conv_std_logic_vector(-571,14),
		conv_std_logic_vector(-565,14),
		conv_std_logic_vector(-558,14),
		conv_std_logic_vector(-552,14),
		conv_std_logic_vector(-546,14),
		conv_std_logic_vector(-539,14),
		conv_std_logic_vector(-533,14),
		conv_std_logic_vector(-527,14),
		conv_std_logic_vector(-521,14),
		conv_std_logic_vector(-514,14),
		conv_std_logic_vector(-508,14),
		conv_std_logic_vector(-502,14),
		conv_std_logic_vector(-496,14),
		conv_std_logic_vector(-489,14),
		conv_std_logic_vector(-483,14),
		conv_std_logic_vector(-477,14),
		conv_std_logic_vector(-470,14),
		conv_std_logic_vector(-464,14),
		conv_std_logic_vector(-458,14),
		conv_std_logic_vector(-452,14),
		conv_std_logic_vector(-445,14),
		conv_std_logic_vector(-439,14),
		conv_std_logic_vector(-433,14),
		conv_std_logic_vector(-427,14),
		conv_std_logic_vector(-420,14),
		conv_std_logic_vector(-414,14),
		conv_std_logic_vector(-408,14),
		conv_std_logic_vector(-401,14),
		conv_std_logic_vector(-395,14),
		conv_std_logic_vector(-389,14),
		conv_std_logic_vector(-383,14),
		conv_std_logic_vector(-376,14),
		conv_std_logic_vector(-370,14),
		conv_std_logic_vector(-364,14),
		conv_std_logic_vector(-358,14),
		conv_std_logic_vector(-351,14),
		conv_std_logic_vector(-345,14),
		conv_std_logic_vector(-339,14),
		conv_std_logic_vector(-332,14),
		conv_std_logic_vector(-326,14),
		conv_std_logic_vector(-320,14),
		conv_std_logic_vector(-314,14),
		conv_std_logic_vector(-307,14),
		conv_std_logic_vector(-301,14),
		conv_std_logic_vector(-295,14),
		conv_std_logic_vector(-288,14),
		conv_std_logic_vector(-282,14),
		conv_std_logic_vector(-276,14),
		conv_std_logic_vector(-270,14),
		conv_std_logic_vector(-263,14),
		conv_std_logic_vector(-257,14),
		conv_std_logic_vector(-251,14),
		conv_std_logic_vector(-245,14),
		conv_std_logic_vector(-238,14),
		conv_std_logic_vector(-232,14),
		conv_std_logic_vector(-226,14),
		conv_std_logic_vector(-219,14),
		conv_std_logic_vector(-213,14),
		conv_std_logic_vector(-207,14),
		conv_std_logic_vector(-201,14),
		conv_std_logic_vector(-194,14),
		conv_std_logic_vector(-188,14),
		conv_std_logic_vector(-182,14),
		conv_std_logic_vector(-175,14),
		conv_std_logic_vector(-169,14),
		conv_std_logic_vector(-163,14),
		conv_std_logic_vector(-157,14),
		conv_std_logic_vector(-150,14),
		conv_std_logic_vector(-144,14),
		conv_std_logic_vector(-138,14),
		conv_std_logic_vector(-131,14),
		conv_std_logic_vector(-125,14),
		conv_std_logic_vector(-119,14),
		conv_std_logic_vector(-113,14),
		conv_std_logic_vector(-106,14),
		conv_std_logic_vector(-100,14),
		conv_std_logic_vector(-94,14),
		conv_std_logic_vector(-87,14),
		conv_std_logic_vector(-81,14),
		conv_std_logic_vector(-75,14),
		conv_std_logic_vector(-69,14),
		conv_std_logic_vector(-62,14),
		conv_std_logic_vector(-56,14),
		conv_std_logic_vector(-50,14),
		conv_std_logic_vector(-43,14),
		conv_std_logic_vector(-37,14),
		conv_std_logic_vector(-31,14),
		conv_std_logic_vector(-25,14),
		conv_std_logic_vector(-18,14),
		conv_std_logic_vector(-12,14),
		conv_std_logic_vector(-6,14));
	signal sdata_out1:	std_logic_vector(27 downto 0);
	signal sdata_out2:	std_logic_vector(27 downto 0);
begin
	
	sdata_out1 <= rom(conv_integer(address1)) * amplitude1;
	data_out1 <= sdata_out1(27 downto 14);
	
	sdata_out2 <= rom(conv_integer(address2)) * amplitude2;
	data_out2 <= sdata_out2(27 downto 14);
	
end;

-- SubModule: sin_counter --

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity sin_counter is
port(
	reset:	in	std_logic;
	clk:	in	std_logic;
	phase_inc:	in	std_logic_vector(12 downto 0);
	Q:		out	std_logic_vector(12 downto 0));
end;

architecture one of sin_counter is
	signal count:	std_logic_vector(12 downto 0);
begin
	Q <= count;
	process(reset,clk)begin
		if(reset = '1')then
			count <= (others => '0');
		elsif(clk 'event and clk = '1')then
			if(count > x"1FFF")then
				count <= (others=>'0');
			else
				count <= count + phase_inc;
			end if;
		end if;
	end process;
end;

-- SubModule: sin_Gen_Peripheral_Register --

library ieee;
use ieee.std_logic_1164.all;

entity sin_Gen_Peripheral_Register is
generic(Bits:integer:=32);
port(
	reset:	in	std_logic;
	clk:	in	std_logic;
	En:		in	std_logic;
	input:	in	std_logic_vector(Bits-1 downto 0);
	output:	out	std_logic_vector(Bits-1 downto 0));
end;

architecture one of sin_Gen_Peripheral_Register is
begin
	process(reset,clk)begin
		if(reset = '1')then
			output <= (others=>'0');
		elsif(clk 'event and clk = '1')then
			if(En = '1')then
				output <= input;
			end if;
		end if;
	end process;
end;